module apb_slave_memory (pclk,
    penable,
    pready,
    prst_n,
    pselx,
    pslverr,
    pwrite,
    paddr,
    prdata,
    pwdata,
    temp);
 input pclk;
 input penable;
 output pready;
 input prst_n;
 input pselx;
 output pslverr;
 input pwrite;
 input [31:0] paddr;
 output [31:0] prdata;
 input [31:0] pwdata;
 output [31:0] temp;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire clknet_leaf_0_pclk;
 wire clknet_leaf_1_pclk;
 wire clknet_leaf_2_pclk;
 wire clknet_leaf_3_pclk;
 wire clknet_leaf_4_pclk;
 wire clknet_leaf_5_pclk;
 wire clknet_leaf_6_pclk;
 wire clknet_leaf_7_pclk;
 wire clknet_leaf_8_pclk;
 wire clknet_leaf_9_pclk;
 wire clknet_leaf_10_pclk;
 wire clknet_leaf_11_pclk;
 wire clknet_leaf_12_pclk;
 wire clknet_leaf_13_pclk;
 wire clknet_leaf_14_pclk;
 wire clknet_leaf_15_pclk;
 wire clknet_leaf_16_pclk;
 wire clknet_leaf_17_pclk;
 wire clknet_leaf_18_pclk;
 wire clknet_leaf_19_pclk;
 wire clknet_leaf_20_pclk;
 wire clknet_leaf_21_pclk;
 wire clknet_leaf_22_pclk;
 wire clknet_leaf_23_pclk;
 wire clknet_leaf_24_pclk;
 wire clknet_leaf_25_pclk;
 wire clknet_leaf_26_pclk;
 wire clknet_leaf_27_pclk;
 wire clknet_leaf_28_pclk;
 wire clknet_leaf_29_pclk;
 wire clknet_leaf_30_pclk;
 wire clknet_leaf_31_pclk;
 wire clknet_leaf_32_pclk;
 wire clknet_leaf_33_pclk;
 wire clknet_leaf_34_pclk;
 wire clknet_leaf_35_pclk;
 wire clknet_0_pclk;
 wire clknet_2_0__leaf_pclk;
 wire clknet_2_1__leaf_pclk;
 wire clknet_2_2__leaf_pclk;
 wire clknet_2_3__leaf_pclk;
 wire net71;
 wire [0:0] _2855_;
 wire [31:0] \mem[0] ;
 wire [31:0] \mem[10] ;
 wire [31:0] \mem[11] ;
 wire [31:0] \mem[12] ;
 wire [31:0] \mem[13] ;
 wire [31:0] \mem[14] ;
 wire [31:0] \mem[15] ;
 wire [31:0] \mem[16] ;
 wire [31:0] \mem[17] ;
 wire [31:0] \mem[18] ;
 wire [31:0] \mem[19] ;
 wire [31:0] \mem[1] ;
 wire [31:0] \mem[20] ;
 wire [31:0] \mem[21] ;
 wire [31:0] \mem[22] ;
 wire [31:0] \mem[23] ;
 wire [31:0] \mem[24] ;
 wire [31:0] \mem[25] ;
 wire [31:0] \mem[26] ;
 wire [31:0] \mem[27] ;
 wire [31:0] \mem[28] ;
 wire [31:0] \mem[29] ;
 wire [31:0] \mem[2] ;
 wire [31:0] \mem[30] ;
 wire [31:0] \mem[31] ;
 wire [31:0] \mem[3] ;
 wire [31:0] \mem[4] ;
 wire [31:0] \mem[5] ;
 wire [31:0] \mem[6] ;
 wire [31:0] \mem[7] ;
 wire [31:0] \mem[8] ;
 wire [31:0] \mem[9] ;
 wire [1:0] next_state;
 wire [1:0] present_state;

 MUX2_X1 _2856_ (.A(pwdata[18]),
    .B(\mem[31] [18]),
    .S(_1102_),
    .Z(_0148_));
 MUX2_X1 _2857_ (.A(pwdata[19]),
    .B(\mem[31] [19]),
    .S(_1102_),
    .Z(_0149_));
 MUX2_X1 _2858_ (.A(pwdata[20]),
    .B(\mem[31] [20]),
    .S(_1102_),
    .Z(_0150_));
 MUX2_X1 _2859_ (.A(pwdata[21]),
    .B(\mem[31] [21]),
    .S(_1102_),
    .Z(_0151_));
 MUX2_X1 _2860_ (.A(pwdata[22]),
    .B(\mem[31] [22]),
    .S(_1102_),
    .Z(_0152_));
 MUX2_X1 _2861_ (.A(pwdata[23]),
    .B(\mem[31] [23]),
    .S(_1102_),
    .Z(_0153_));
 MUX2_X1 _2862_ (.A(pwdata[24]),
    .B(\mem[31] [24]),
    .S(_1102_),
    .Z(_0154_));
 MUX2_X1 _2863_ (.A(pwdata[25]),
    .B(\mem[31] [25]),
    .S(_1102_),
    .Z(_0155_));
 MUX2_X1 _2864_ (.A(pwdata[26]),
    .B(\mem[31] [26]),
    .S(_1102_),
    .Z(_0156_));
 MUX2_X1 _2865_ (.A(pwdata[27]),
    .B(\mem[31] [27]),
    .S(_1102_),
    .Z(_0157_));
 MUX2_X1 _2866_ (.A(pwdata[28]),
    .B(\mem[31] [28]),
    .S(_1102_),
    .Z(_0158_));
 MUX2_X1 _2867_ (.A(pwdata[29]),
    .B(\mem[31] [29]),
    .S(_1102_),
    .Z(_0159_));
 MUX2_X1 _2868_ (.A(pwdata[30]),
    .B(\mem[31] [30]),
    .S(_1102_),
    .Z(_0160_));
 MUX2_X1 _2869_ (.A(pwdata[31]),
    .B(\mem[31] [31]),
    .S(_1102_),
    .Z(_0161_));
 NOR4_X4 _2870_ (.A1(_1069_),
    .A2(paddr[1]),
    .A3(_1073_),
    .A4(_1098_),
    .ZN(_1103_));
 NAND2_X4 _2871_ (.A1(_1090_),
    .A2(net69),
    .ZN(_1104_));
 MUX2_X1 _2872_ (.A(pwdata[0]),
    .B(\mem[17] [0]),
    .S(_1104_),
    .Z(_0162_));
 MUX2_X1 _2873_ (.A(pwdata[1]),
    .B(\mem[17] [1]),
    .S(_1104_),
    .Z(_0163_));
 MUX2_X1 _2874_ (.A(pwdata[2]),
    .B(\mem[17] [2]),
    .S(_1104_),
    .Z(_0164_));
 MUX2_X1 _2875_ (.A(pwdata[3]),
    .B(\mem[17] [3]),
    .S(_1104_),
    .Z(_0165_));
 MUX2_X1 _2876_ (.A(pwdata[4]),
    .B(\mem[17] [4]),
    .S(_1104_),
    .Z(_0166_));
 MUX2_X1 _2877_ (.A(pwdata[5]),
    .B(\mem[17] [5]),
    .S(_1104_),
    .Z(_0167_));
 MUX2_X1 _2878_ (.A(pwdata[6]),
    .B(\mem[17] [6]),
    .S(_1104_),
    .Z(_0168_));
 MUX2_X1 _2879_ (.A(pwdata[7]),
    .B(\mem[17] [7]),
    .S(_1104_),
    .Z(_0169_));
 MUX2_X1 _2880_ (.A(pwdata[8]),
    .B(\mem[17] [8]),
    .S(_1104_),
    .Z(_0170_));
 MUX2_X1 _2881_ (.A(pwdata[9]),
    .B(\mem[17] [9]),
    .S(_1104_),
    .Z(_0171_));
 MUX2_X1 _2882_ (.A(pwdata[10]),
    .B(\mem[17] [10]),
    .S(_1104_),
    .Z(_0172_));
 MUX2_X1 _2883_ (.A(pwdata[11]),
    .B(\mem[17] [11]),
    .S(_1104_),
    .Z(_0173_));
 MUX2_X1 _2884_ (.A(pwdata[12]),
    .B(\mem[17] [12]),
    .S(_1104_),
    .Z(_0174_));
 MUX2_X1 _2885_ (.A(pwdata[13]),
    .B(\mem[17] [13]),
    .S(_1104_),
    .Z(_0175_));
 MUX2_X1 _2886_ (.A(pwdata[14]),
    .B(\mem[17] [14]),
    .S(_1104_),
    .Z(_0176_));
 MUX2_X1 _2887_ (.A(pwdata[15]),
    .B(\mem[17] [15]),
    .S(_1104_),
    .Z(_0177_));
 MUX2_X1 _2888_ (.A(pwdata[16]),
    .B(\mem[17] [16]),
    .S(_1104_),
    .Z(_0178_));
 MUX2_X1 _2889_ (.A(pwdata[17]),
    .B(\mem[17] [17]),
    .S(_1104_),
    .Z(_0179_));
 MUX2_X1 _2890_ (.A(pwdata[18]),
    .B(\mem[17] [18]),
    .S(_1104_),
    .Z(_0180_));
 MUX2_X1 _2891_ (.A(pwdata[19]),
    .B(\mem[17] [19]),
    .S(_1104_),
    .Z(_0181_));
 MUX2_X1 _2892_ (.A(pwdata[20]),
    .B(\mem[17] [20]),
    .S(_1104_),
    .Z(_0182_));
 MUX2_X1 _2893_ (.A(pwdata[21]),
    .B(\mem[17] [21]),
    .S(_1104_),
    .Z(_0183_));
 MUX2_X1 _2894_ (.A(pwdata[22]),
    .B(\mem[17] [22]),
    .S(_1104_),
    .Z(_0184_));
 MUX2_X1 _2895_ (.A(pwdata[23]),
    .B(\mem[17] [23]),
    .S(_1104_),
    .Z(_0185_));
 MUX2_X1 _2896_ (.A(pwdata[24]),
    .B(\mem[17] [24]),
    .S(_1104_),
    .Z(_0186_));
 MUX2_X1 _2897_ (.A(pwdata[25]),
    .B(\mem[17] [25]),
    .S(_1104_),
    .Z(_0187_));
 MUX2_X1 _2898_ (.A(pwdata[26]),
    .B(\mem[17] [26]),
    .S(_1104_),
    .Z(_0188_));
 MUX2_X1 _2899_ (.A(pwdata[27]),
    .B(\mem[17] [27]),
    .S(_1104_),
    .Z(_0189_));
 MUX2_X1 _2900_ (.A(pwdata[28]),
    .B(\mem[17] [28]),
    .S(_1104_),
    .Z(_0190_));
 MUX2_X1 _2901_ (.A(pwdata[29]),
    .B(\mem[17] [29]),
    .S(_1104_),
    .Z(_0191_));
 MUX2_X1 _2902_ (.A(pwdata[30]),
    .B(\mem[17] [30]),
    .S(_1104_),
    .Z(_0192_));
 MUX2_X1 _2903_ (.A(pwdata[31]),
    .B(\mem[17] [31]),
    .S(_1104_),
    .Z(_0193_));
 NOR4_X4 _2904_ (.A1(_1069_),
    .A2(_1070_),
    .A3(paddr[2]),
    .A4(_1092_),
    .ZN(_1105_));
 NAND2_X4 _2905_ (.A1(_1090_),
    .A2(net67),
    .ZN(_1106_));
 MUX2_X1 _2906_ (.A(pwdata[0]),
    .B(\mem[27] [0]),
    .S(_1106_),
    .Z(_0194_));
 MUX2_X1 _2907_ (.A(pwdata[1]),
    .B(\mem[27] [1]),
    .S(_1106_),
    .Z(_0195_));
 MUX2_X1 _2908_ (.A(pwdata[2]),
    .B(\mem[27] [2]),
    .S(_1106_),
    .Z(_0196_));
 MUX2_X1 _2909_ (.A(pwdata[3]),
    .B(\mem[27] [3]),
    .S(_1106_),
    .Z(_0197_));
 MUX2_X1 _2910_ (.A(pwdata[4]),
    .B(\mem[27] [4]),
    .S(_1106_),
    .Z(_0198_));
 MUX2_X1 _2911_ (.A(pwdata[5]),
    .B(\mem[27] [5]),
    .S(_1106_),
    .Z(_0199_));
 MUX2_X1 _2912_ (.A(pwdata[6]),
    .B(\mem[27] [6]),
    .S(_1106_),
    .Z(_0200_));
 MUX2_X1 _2913_ (.A(pwdata[7]),
    .B(\mem[27] [7]),
    .S(_1106_),
    .Z(_0201_));
 MUX2_X1 _2914_ (.A(pwdata[8]),
    .B(\mem[27] [8]),
    .S(_1106_),
    .Z(_0202_));
 MUX2_X1 _2915_ (.A(pwdata[9]),
    .B(\mem[27] [9]),
    .S(_1106_),
    .Z(_0203_));
 MUX2_X1 _2916_ (.A(pwdata[10]),
    .B(\mem[27] [10]),
    .S(_1106_),
    .Z(_0204_));
 MUX2_X1 _2917_ (.A(pwdata[11]),
    .B(\mem[27] [11]),
    .S(_1106_),
    .Z(_0205_));
 MUX2_X1 _2918_ (.A(pwdata[12]),
    .B(\mem[27] [12]),
    .S(_1106_),
    .Z(_0206_));
 MUX2_X1 _2919_ (.A(pwdata[13]),
    .B(\mem[27] [13]),
    .S(_1106_),
    .Z(_0207_));
 MUX2_X1 _2920_ (.A(pwdata[14]),
    .B(\mem[27] [14]),
    .S(_1106_),
    .Z(_0208_));
 MUX2_X1 _2921_ (.A(pwdata[15]),
    .B(\mem[27] [15]),
    .S(_1106_),
    .Z(_0209_));
 MUX2_X1 _2922_ (.A(pwdata[16]),
    .B(\mem[27] [16]),
    .S(_1106_),
    .Z(_0210_));
 MUX2_X1 _2923_ (.A(pwdata[17]),
    .B(\mem[27] [17]),
    .S(_1106_),
    .Z(_0211_));
 MUX2_X1 _2924_ (.A(pwdata[18]),
    .B(\mem[27] [18]),
    .S(_1106_),
    .Z(_0212_));
 MUX2_X1 _2925_ (.A(pwdata[19]),
    .B(\mem[27] [19]),
    .S(_1106_),
    .Z(_0213_));
 MUX2_X1 _2926_ (.A(pwdata[20]),
    .B(\mem[27] [20]),
    .S(_1106_),
    .Z(_0214_));
 MUX2_X1 _2927_ (.A(pwdata[21]),
    .B(\mem[27] [21]),
    .S(_1106_),
    .Z(_0215_));
 MUX2_X1 _2928_ (.A(pwdata[22]),
    .B(\mem[27] [22]),
    .S(_1106_),
    .Z(_0216_));
 MUX2_X1 _2929_ (.A(pwdata[23]),
    .B(\mem[27] [23]),
    .S(_1106_),
    .Z(_0217_));
 MUX2_X1 _2930_ (.A(pwdata[24]),
    .B(\mem[27] [24]),
    .S(_1106_),
    .Z(_0218_));
 MUX2_X1 _2931_ (.A(pwdata[25]),
    .B(\mem[27] [25]),
    .S(_1106_),
    .Z(_0219_));
 MUX2_X1 _2932_ (.A(pwdata[26]),
    .B(\mem[27] [26]),
    .S(_1106_),
    .Z(_0220_));
 MUX2_X1 _2933_ (.A(pwdata[27]),
    .B(\mem[27] [27]),
    .S(_1106_),
    .Z(_0221_));
 MUX2_X1 _2934_ (.A(pwdata[28]),
    .B(\mem[27] [28]),
    .S(_1106_),
    .Z(_0222_));
 MUX2_X1 _2935_ (.A(pwdata[29]),
    .B(\mem[27] [29]),
    .S(_1106_),
    .Z(_0223_));
 MUX2_X1 _2936_ (.A(pwdata[30]),
    .B(\mem[27] [30]),
    .S(_1106_),
    .Z(_0224_));
 MUX2_X1 _2937_ (.A(pwdata[31]),
    .B(\mem[27] [31]),
    .S(_1106_),
    .Z(_0225_));
 NOR4_X4 _2938_ (.A1(_1069_),
    .A2(_1072_),
    .A3(paddr[0]),
    .A4(_1098_),
    .ZN(_1107_));
 NAND2_X4 _2939_ (.A1(net2),
    .A2(net65),
    .ZN(_1108_));
 MUX2_X1 _2940_ (.A(pwdata[0]),
    .B(\mem[18] [0]),
    .S(_1108_),
    .Z(_0226_));
 MUX2_X1 _2941_ (.A(pwdata[1]),
    .B(\mem[18] [1]),
    .S(_1108_),
    .Z(_0227_));
 MUX2_X1 _2942_ (.A(pwdata[2]),
    .B(\mem[18] [2]),
    .S(_1108_),
    .Z(_0228_));
 MUX2_X1 _2943_ (.A(pwdata[3]),
    .B(\mem[18] [3]),
    .S(_1108_),
    .Z(_0229_));
 MUX2_X1 _2944_ (.A(pwdata[4]),
    .B(\mem[18] [4]),
    .S(_1108_),
    .Z(_0230_));
 MUX2_X1 _2945_ (.A(pwdata[5]),
    .B(\mem[18] [5]),
    .S(_1108_),
    .Z(_0231_));
 MUX2_X1 _2946_ (.A(pwdata[6]),
    .B(\mem[18] [6]),
    .S(_1108_),
    .Z(_0232_));
 MUX2_X1 _2947_ (.A(pwdata[7]),
    .B(\mem[18] [7]),
    .S(_1108_),
    .Z(_0233_));
 MUX2_X1 _2948_ (.A(pwdata[8]),
    .B(\mem[18] [8]),
    .S(_1108_),
    .Z(_0234_));
 MUX2_X1 _2949_ (.A(pwdata[9]),
    .B(\mem[18] [9]),
    .S(_1108_),
    .Z(_0235_));
 MUX2_X1 _2950_ (.A(pwdata[10]),
    .B(\mem[18] [10]),
    .S(_1108_),
    .Z(_0236_));
 MUX2_X1 _2951_ (.A(pwdata[11]),
    .B(\mem[18] [11]),
    .S(_1108_),
    .Z(_0237_));
 MUX2_X1 _2952_ (.A(pwdata[12]),
    .B(\mem[18] [12]),
    .S(_1108_),
    .Z(_0238_));
 MUX2_X1 _2953_ (.A(pwdata[13]),
    .B(\mem[18] [13]),
    .S(_1108_),
    .Z(_0239_));
 MUX2_X1 _2954_ (.A(pwdata[14]),
    .B(\mem[18] [14]),
    .S(_1108_),
    .Z(_0240_));
 MUX2_X1 _2955_ (.A(pwdata[15]),
    .B(\mem[18] [15]),
    .S(_1108_),
    .Z(_0241_));
 MUX2_X1 _2956_ (.A(pwdata[16]),
    .B(\mem[18] [16]),
    .S(_1108_),
    .Z(_0242_));
 MUX2_X1 _2957_ (.A(pwdata[17]),
    .B(\mem[18] [17]),
    .S(_1108_),
    .Z(_0243_));
 MUX2_X1 _2958_ (.A(pwdata[18]),
    .B(\mem[18] [18]),
    .S(_1108_),
    .Z(_0244_));
 MUX2_X1 _2959_ (.A(pwdata[19]),
    .B(\mem[18] [19]),
    .S(_1108_),
    .Z(_0245_));
 MUX2_X1 _2960_ (.A(pwdata[20]),
    .B(\mem[18] [20]),
    .S(_1108_),
    .Z(_0246_));
 MUX2_X1 _2961_ (.A(pwdata[21]),
    .B(\mem[18] [21]),
    .S(_1108_),
    .Z(_0247_));
 MUX2_X1 _2962_ (.A(pwdata[22]),
    .B(\mem[18] [22]),
    .S(_1108_),
    .Z(_0248_));
 MUX2_X1 _2963_ (.A(pwdata[23]),
    .B(\mem[18] [23]),
    .S(_1108_),
    .Z(_0249_));
 MUX2_X1 _2964_ (.A(pwdata[24]),
    .B(\mem[18] [24]),
    .S(_1108_),
    .Z(_0250_));
 MUX2_X1 _2965_ (.A(pwdata[25]),
    .B(\mem[18] [25]),
    .S(_1108_),
    .Z(_0251_));
 MUX2_X1 _2966_ (.A(pwdata[26]),
    .B(\mem[18] [26]),
    .S(_1108_),
    .Z(_0252_));
 MUX2_X1 _2967_ (.A(pwdata[27]),
    .B(\mem[18] [27]),
    .S(_1108_),
    .Z(_0253_));
 MUX2_X1 _2968_ (.A(pwdata[28]),
    .B(\mem[18] [28]),
    .S(_1108_),
    .Z(_0254_));
 MUX2_X1 _2969_ (.A(pwdata[29]),
    .B(\mem[18] [29]),
    .S(_1108_),
    .Z(_0255_));
 MUX2_X1 _2970_ (.A(pwdata[30]),
    .B(\mem[18] [30]),
    .S(_1108_),
    .Z(_0256_));
 MUX2_X1 _2971_ (.A(pwdata[31]),
    .B(\mem[18] [31]),
    .S(_1108_),
    .Z(_0257_));
 NOR3_X4 _2972_ (.A1(_1069_),
    .A2(_1075_),
    .A3(_1076_),
    .ZN(_1109_));
 NAND2_X4 _2973_ (.A1(net2),
    .A2(net62),
    .ZN(_1110_));
 MUX2_X1 _2974_ (.A(pwdata[0]),
    .B(\mem[28] [0]),
    .S(_1110_),
    .Z(_0258_));
 MUX2_X1 _2975_ (.A(pwdata[1]),
    .B(\mem[28] [1]),
    .S(_1110_),
    .Z(_0259_));
 MUX2_X1 _2976_ (.A(pwdata[2]),
    .B(\mem[28] [2]),
    .S(_1110_),
    .Z(_0260_));
 MUX2_X1 _2977_ (.A(pwdata[3]),
    .B(\mem[28] [3]),
    .S(_1110_),
    .Z(_0261_));
 MUX2_X1 _2978_ (.A(pwdata[4]),
    .B(\mem[28] [4]),
    .S(_1110_),
    .Z(_0262_));
 MUX2_X1 _2979_ (.A(pwdata[5]),
    .B(\mem[28] [5]),
    .S(_1110_),
    .Z(_0263_));
 MUX2_X1 _2980_ (.A(pwdata[6]),
    .B(\mem[28] [6]),
    .S(_1110_),
    .Z(_0264_));
 MUX2_X1 _2981_ (.A(pwdata[7]),
    .B(\mem[28] [7]),
    .S(_1110_),
    .Z(_0265_));
 MUX2_X1 _2982_ (.A(pwdata[8]),
    .B(\mem[28] [8]),
    .S(_1110_),
    .Z(_0266_));
 MUX2_X1 _2983_ (.A(pwdata[9]),
    .B(\mem[28] [9]),
    .S(_1110_),
    .Z(_0267_));
 MUX2_X1 _2984_ (.A(pwdata[10]),
    .B(\mem[28] [10]),
    .S(_1110_),
    .Z(_0268_));
 MUX2_X1 _2985_ (.A(pwdata[11]),
    .B(\mem[28] [11]),
    .S(_1110_),
    .Z(_0269_));
 MUX2_X1 _2986_ (.A(pwdata[12]),
    .B(\mem[28] [12]),
    .S(_1110_),
    .Z(_0270_));
 MUX2_X1 _2987_ (.A(pwdata[13]),
    .B(\mem[28] [13]),
    .S(_1110_),
    .Z(_0271_));
 MUX2_X1 _2988_ (.A(pwdata[14]),
    .B(\mem[28] [14]),
    .S(_1110_),
    .Z(_0272_));
 MUX2_X1 _2989_ (.A(pwdata[15]),
    .B(\mem[28] [15]),
    .S(_1110_),
    .Z(_0273_));
 MUX2_X1 _2990_ (.A(pwdata[16]),
    .B(\mem[28] [16]),
    .S(_1110_),
    .Z(_0274_));
 MUX2_X1 _2991_ (.A(pwdata[17]),
    .B(\mem[28] [17]),
    .S(_1110_),
    .Z(_0275_));
 MUX2_X1 _2992_ (.A(pwdata[18]),
    .B(\mem[28] [18]),
    .S(_1110_),
    .Z(_0276_));
 MUX2_X1 _2993_ (.A(pwdata[19]),
    .B(\mem[28] [19]),
    .S(_1110_),
    .Z(_0277_));
 MUX2_X1 _2994_ (.A(pwdata[20]),
    .B(\mem[28] [20]),
    .S(_1110_),
    .Z(_0278_));
 MUX2_X1 _2995_ (.A(pwdata[21]),
    .B(\mem[28] [21]),
    .S(_1110_),
    .Z(_0279_));
 MUX2_X1 _2996_ (.A(pwdata[22]),
    .B(\mem[28] [22]),
    .S(_1110_),
    .Z(_0280_));
 MUX2_X1 _2997_ (.A(pwdata[23]),
    .B(\mem[28] [23]),
    .S(_1110_),
    .Z(_0281_));
 MUX2_X1 _2998_ (.A(pwdata[24]),
    .B(\mem[28] [24]),
    .S(_1110_),
    .Z(_0282_));
 MUX2_X1 _2999_ (.A(pwdata[25]),
    .B(\mem[28] [25]),
    .S(_1110_),
    .Z(_0283_));
 MUX2_X1 _3000_ (.A(pwdata[26]),
    .B(\mem[28] [26]),
    .S(_1110_),
    .Z(_0284_));
 MUX2_X1 _3001_ (.A(pwdata[27]),
    .B(\mem[28] [27]),
    .S(_1110_),
    .Z(_0285_));
 MUX2_X1 _3002_ (.A(pwdata[28]),
    .B(\mem[28] [28]),
    .S(_1110_),
    .Z(_0286_));
 MUX2_X1 _3003_ (.A(pwdata[29]),
    .B(\mem[28] [29]),
    .S(_1110_),
    .Z(_0287_));
 MUX2_X1 _3004_ (.A(pwdata[30]),
    .B(\mem[28] [30]),
    .S(_1110_),
    .Z(_0288_));
 MUX2_X1 _3005_ (.A(pwdata[31]),
    .B(\mem[28] [31]),
    .S(_1110_),
    .Z(_0289_));
 NOR3_X4 _3006_ (.A1(_1069_),
    .A2(_1092_),
    .A3(_1098_),
    .ZN(_1111_));
 NAND2_X4 _3007_ (.A1(net2),
    .A2(net59),
    .ZN(_1112_));
 MUX2_X1 _3008_ (.A(pwdata[0]),
    .B(\mem[19] [0]),
    .S(_1112_),
    .Z(_0290_));
 MUX2_X1 _3009_ (.A(pwdata[1]),
    .B(\mem[19] [1]),
    .S(_1112_),
    .Z(_0291_));
 MUX2_X1 _3010_ (.A(pwdata[2]),
    .B(\mem[19] [2]),
    .S(_1112_),
    .Z(_0292_));
 MUX2_X1 _3011_ (.A(pwdata[3]),
    .B(\mem[19] [3]),
    .S(_1112_),
    .Z(_0293_));
 MUX2_X1 _3012_ (.A(pwdata[4]),
    .B(\mem[19] [4]),
    .S(_1112_),
    .Z(_0294_));
 MUX2_X1 _3013_ (.A(pwdata[5]),
    .B(\mem[19] [5]),
    .S(_1112_),
    .Z(_0295_));
 MUX2_X1 _3014_ (.A(pwdata[6]),
    .B(\mem[19] [6]),
    .S(_1112_),
    .Z(_0296_));
 MUX2_X1 _3015_ (.A(pwdata[7]),
    .B(\mem[19] [7]),
    .S(_1112_),
    .Z(_0297_));
 MUX2_X1 _3016_ (.A(pwdata[8]),
    .B(\mem[19] [8]),
    .S(_1112_),
    .Z(_0298_));
 MUX2_X1 _3017_ (.A(pwdata[9]),
    .B(\mem[19] [9]),
    .S(_1112_),
    .Z(_0299_));
 MUX2_X1 _3018_ (.A(pwdata[10]),
    .B(\mem[19] [10]),
    .S(_1112_),
    .Z(_0300_));
 MUX2_X1 _3019_ (.A(pwdata[11]),
    .B(\mem[19] [11]),
    .S(_1112_),
    .Z(_0301_));
 MUX2_X1 _3020_ (.A(pwdata[12]),
    .B(\mem[19] [12]),
    .S(_1112_),
    .Z(_0302_));
 MUX2_X1 _3021_ (.A(pwdata[13]),
    .B(\mem[19] [13]),
    .S(_1112_),
    .Z(_0303_));
 MUX2_X1 _3022_ (.A(pwdata[14]),
    .B(\mem[19] [14]),
    .S(_1112_),
    .Z(_0304_));
 MUX2_X1 _3023_ (.A(pwdata[15]),
    .B(\mem[19] [15]),
    .S(_1112_),
    .Z(_0305_));
 MUX2_X1 _3024_ (.A(pwdata[16]),
    .B(\mem[19] [16]),
    .S(_1112_),
    .Z(_0306_));
 MUX2_X1 _3025_ (.A(pwdata[17]),
    .B(\mem[19] [17]),
    .S(_1112_),
    .Z(_0307_));
 MUX2_X1 _3026_ (.A(pwdata[18]),
    .B(\mem[19] [18]),
    .S(_1112_),
    .Z(_0308_));
 MUX2_X1 _3027_ (.A(pwdata[19]),
    .B(\mem[19] [19]),
    .S(_1112_),
    .Z(_0309_));
 MUX2_X1 _3028_ (.A(pwdata[20]),
    .B(\mem[19] [20]),
    .S(_1112_),
    .Z(_0310_));
 MUX2_X1 _3029_ (.A(pwdata[21]),
    .B(\mem[19] [21]),
    .S(_1112_),
    .Z(_0311_));
 MUX2_X1 _3030_ (.A(pwdata[22]),
    .B(\mem[19] [22]),
    .S(_1112_),
    .Z(_0312_));
 MUX2_X1 _3031_ (.A(pwdata[23]),
    .B(\mem[19] [23]),
    .S(_1112_),
    .Z(_0313_));
 MUX2_X1 _3032_ (.A(pwdata[24]),
    .B(\mem[19] [24]),
    .S(_1112_),
    .Z(_0314_));
 MUX2_X1 _3033_ (.A(pwdata[25]),
    .B(\mem[19] [25]),
    .S(_1112_),
    .Z(_0315_));
 MUX2_X1 _3034_ (.A(pwdata[26]),
    .B(\mem[19] [26]),
    .S(_1112_),
    .Z(_0316_));
 MUX2_X1 _3035_ (.A(pwdata[27]),
    .B(\mem[19] [27]),
    .S(_1112_),
    .Z(_0317_));
 MUX2_X1 _3036_ (.A(pwdata[28]),
    .B(\mem[19] [28]),
    .S(_1112_),
    .Z(_0318_));
 MUX2_X1 _3037_ (.A(pwdata[29]),
    .B(\mem[19] [29]),
    .S(_1112_),
    .Z(_0319_));
 MUX2_X1 _3038_ (.A(pwdata[30]),
    .B(\mem[19] [30]),
    .S(_1112_),
    .Z(_0320_));
 MUX2_X1 _3039_ (.A(pwdata[31]),
    .B(\mem[19] [31]),
    .S(_1112_),
    .Z(_0321_));
 NOR4_X4 _3040_ (.A1(_1069_),
    .A2(_1070_),
    .A3(paddr[2]),
    .A4(_1076_),
    .ZN(_1113_));
 NAND2_X4 _3041_ (.A1(net2),
    .A2(net58),
    .ZN(_1114_));
 MUX2_X1 _3042_ (.A(pwdata[0]),
    .B(\mem[24] [0]),
    .S(_1114_),
    .Z(_0322_));
 MUX2_X1 _3043_ (.A(pwdata[1]),
    .B(\mem[24] [1]),
    .S(_1114_),
    .Z(_0323_));
 MUX2_X1 _3044_ (.A(pwdata[2]),
    .B(\mem[24] [2]),
    .S(_1114_),
    .Z(_0324_));
 MUX2_X1 _3045_ (.A(pwdata[3]),
    .B(\mem[24] [3]),
    .S(_1114_),
    .Z(_0325_));
 MUX2_X1 _3046_ (.A(pwdata[4]),
    .B(\mem[24] [4]),
    .S(_1114_),
    .Z(_0326_));
 MUX2_X1 _3047_ (.A(pwdata[5]),
    .B(\mem[24] [5]),
    .S(_1114_),
    .Z(_0327_));
 MUX2_X1 _3048_ (.A(pwdata[6]),
    .B(\mem[24] [6]),
    .S(_1114_),
    .Z(_0328_));
 MUX2_X1 _3049_ (.A(pwdata[7]),
    .B(\mem[24] [7]),
    .S(_1114_),
    .Z(_0329_));
 MUX2_X1 _3050_ (.A(pwdata[8]),
    .B(\mem[24] [8]),
    .S(_1114_),
    .Z(_0330_));
 MUX2_X1 _3051_ (.A(pwdata[9]),
    .B(\mem[24] [9]),
    .S(_1114_),
    .Z(_0331_));
 MUX2_X1 _3052_ (.A(pwdata[10]),
    .B(\mem[24] [10]),
    .S(_1114_),
    .Z(_0332_));
 MUX2_X1 _3053_ (.A(pwdata[11]),
    .B(\mem[24] [11]),
    .S(_1114_),
    .Z(_0333_));
 MUX2_X1 _3054_ (.A(pwdata[12]),
    .B(\mem[24] [12]),
    .S(_1114_),
    .Z(_0334_));
 MUX2_X1 _3055_ (.A(pwdata[13]),
    .B(\mem[24] [13]),
    .S(_1114_),
    .Z(_0335_));
 MUX2_X1 _3056_ (.A(pwdata[14]),
    .B(\mem[24] [14]),
    .S(_1114_),
    .Z(_0336_));
 MUX2_X1 _3057_ (.A(pwdata[15]),
    .B(\mem[24] [15]),
    .S(_1114_),
    .Z(_0337_));
 MUX2_X1 _3058_ (.A(pwdata[16]),
    .B(\mem[24] [16]),
    .S(_1114_),
    .Z(_0338_));
 MUX2_X1 _3059_ (.A(pwdata[17]),
    .B(\mem[24] [17]),
    .S(_1114_),
    .Z(_0339_));
 MUX2_X1 _3060_ (.A(pwdata[18]),
    .B(\mem[24] [18]),
    .S(_1114_),
    .Z(_0340_));
 MUX2_X1 _3061_ (.A(pwdata[19]),
    .B(\mem[24] [19]),
    .S(_1114_),
    .Z(_0341_));
 MUX2_X1 _3062_ (.A(pwdata[20]),
    .B(\mem[24] [20]),
    .S(_1114_),
    .Z(_0342_));
 MUX2_X1 _3063_ (.A(pwdata[21]),
    .B(\mem[24] [21]),
    .S(_1114_),
    .Z(_0343_));
 MUX2_X1 _3064_ (.A(pwdata[22]),
    .B(\mem[24] [22]),
    .S(_1114_),
    .Z(_0344_));
 MUX2_X1 _3065_ (.A(pwdata[23]),
    .B(\mem[24] [23]),
    .S(_1114_),
    .Z(_0345_));
 MUX2_X1 _3066_ (.A(pwdata[24]),
    .B(\mem[24] [24]),
    .S(_1114_),
    .Z(_0346_));
 MUX2_X1 _3067_ (.A(pwdata[25]),
    .B(\mem[24] [25]),
    .S(_1114_),
    .Z(_0347_));
 MUX2_X1 _3068_ (.A(pwdata[26]),
    .B(\mem[24] [26]),
    .S(_1114_),
    .Z(_0348_));
 MUX2_X1 _3069_ (.A(pwdata[27]),
    .B(\mem[24] [27]),
    .S(_1114_),
    .Z(_0349_));
 MUX2_X1 _3070_ (.A(pwdata[28]),
    .B(\mem[24] [28]),
    .S(_1114_),
    .Z(_0350_));
 MUX2_X1 _3071_ (.A(pwdata[29]),
    .B(\mem[24] [29]),
    .S(_1114_),
    .Z(_0351_));
 MUX2_X1 _3072_ (.A(pwdata[30]),
    .B(\mem[24] [30]),
    .S(_1114_),
    .Z(_0352_));
 MUX2_X1 _3073_ (.A(pwdata[31]),
    .B(\mem[24] [31]),
    .S(_1114_),
    .Z(_0353_));
 NOR4_X1 _3074_ (.A1(_1070_),
    .A2(paddr[2]),
    .A3(paddr[1]),
    .A4(_1073_),
    .ZN(_1115_));
 AND2_X2 _3075_ (.A1(_1069_),
    .A2(_1115_),
    .ZN(_1116_));
 NAND2_X4 _3076_ (.A1(net2),
    .A2(net5),
    .ZN(_1117_));
 MUX2_X1 _3077_ (.A(pwdata[0]),
    .B(\mem[9] [0]),
    .S(_1117_),
    .Z(_0354_));
 MUX2_X1 _3078_ (.A(pwdata[1]),
    .B(\mem[9] [1]),
    .S(_1117_),
    .Z(_0355_));
 MUX2_X1 _3079_ (.A(pwdata[2]),
    .B(\mem[9] [2]),
    .S(_1117_),
    .Z(_0356_));
 MUX2_X1 _3080_ (.A(pwdata[3]),
    .B(\mem[9] [3]),
    .S(_1117_),
    .Z(_0357_));
 MUX2_X1 _3081_ (.A(pwdata[4]),
    .B(\mem[9] [4]),
    .S(_1117_),
    .Z(_0358_));
 MUX2_X1 _3082_ (.A(pwdata[5]),
    .B(\mem[9] [5]),
    .S(_1117_),
    .Z(_0359_));
 MUX2_X1 _3083_ (.A(pwdata[6]),
    .B(\mem[9] [6]),
    .S(_1117_),
    .Z(_0360_));
 MUX2_X1 _3084_ (.A(pwdata[7]),
    .B(\mem[9] [7]),
    .S(_1117_),
    .Z(_0361_));
 MUX2_X1 _3085_ (.A(pwdata[8]),
    .B(\mem[9] [8]),
    .S(_1117_),
    .Z(_0362_));
 MUX2_X1 _3086_ (.A(pwdata[9]),
    .B(\mem[9] [9]),
    .S(_1117_),
    .Z(_0363_));
 MUX2_X1 _3087_ (.A(pwdata[10]),
    .B(\mem[9] [10]),
    .S(_1117_),
    .Z(_0364_));
 MUX2_X1 _3088_ (.A(pwdata[11]),
    .B(\mem[9] [11]),
    .S(_1117_),
    .Z(_0365_));
 MUX2_X1 _3089_ (.A(pwdata[12]),
    .B(\mem[9] [12]),
    .S(_1117_),
    .Z(_0366_));
 MUX2_X1 _3090_ (.A(pwdata[13]),
    .B(\mem[9] [13]),
    .S(_1117_),
    .Z(_0367_));
 MUX2_X1 _3091_ (.A(pwdata[14]),
    .B(\mem[9] [14]),
    .S(_1117_),
    .Z(_0368_));
 MUX2_X1 _3092_ (.A(pwdata[15]),
    .B(\mem[9] [15]),
    .S(_1117_),
    .Z(_0369_));
 MUX2_X1 _3093_ (.A(pwdata[16]),
    .B(\mem[9] [16]),
    .S(_1117_),
    .Z(_0370_));
 MUX2_X1 _3094_ (.A(pwdata[17]),
    .B(\mem[9] [17]),
    .S(_1117_),
    .Z(_0371_));
 MUX2_X1 _3095_ (.A(pwdata[18]),
    .B(\mem[9] [18]),
    .S(_1117_),
    .Z(_0372_));
 MUX2_X1 _3096_ (.A(pwdata[19]),
    .B(\mem[9] [19]),
    .S(_1117_),
    .Z(_0373_));
 MUX2_X1 _3097_ (.A(pwdata[20]),
    .B(\mem[9] [20]),
    .S(_1117_),
    .Z(_0374_));
 MUX2_X1 _3098_ (.A(pwdata[21]),
    .B(\mem[9] [21]),
    .S(_1117_),
    .Z(_0375_));
 MUX2_X1 _3099_ (.A(pwdata[22]),
    .B(\mem[9] [22]),
    .S(_1117_),
    .Z(_0376_));
 MUX2_X1 _3100_ (.A(pwdata[23]),
    .B(\mem[9] [23]),
    .S(_1117_),
    .Z(_0377_));
 MUX2_X1 _3101_ (.A(pwdata[24]),
    .B(\mem[9] [24]),
    .S(_1117_),
    .Z(_0378_));
 MUX2_X1 _3102_ (.A(pwdata[25]),
    .B(\mem[9] [25]),
    .S(_1117_),
    .Z(_0379_));
 MUX2_X1 _3103_ (.A(pwdata[26]),
    .B(\mem[9] [26]),
    .S(_1117_),
    .Z(_0380_));
 MUX2_X1 _3104_ (.A(pwdata[27]),
    .B(\mem[9] [27]),
    .S(_1117_),
    .Z(_0381_));
 MUX2_X1 _3105_ (.A(pwdata[28]),
    .B(\mem[9] [28]),
    .S(_1117_),
    .Z(_0382_));
 MUX2_X1 _3106_ (.A(pwdata[29]),
    .B(\mem[9] [29]),
    .S(_1117_),
    .Z(_0383_));
 MUX2_X1 _3107_ (.A(pwdata[30]),
    .B(\mem[9] [30]),
    .S(_1117_),
    .Z(_0384_));
 MUX2_X1 _3108_ (.A(pwdata[31]),
    .B(\mem[9] [31]),
    .S(_1117_),
    .Z(_0385_));
 NOR4_X4 _3109_ (.A1(_1069_),
    .A2(paddr[3]),
    .A3(_1071_),
    .A4(_1076_),
    .ZN(_1118_));
 NAND2_X4 _3110_ (.A1(_1090_),
    .A2(net53),
    .ZN(_1119_));
 MUX2_X1 _3111_ (.A(pwdata[0]),
    .B(\mem[20] [0]),
    .S(_1119_),
    .Z(_0386_));
 MUX2_X1 _3112_ (.A(pwdata[1]),
    .B(\mem[20] [1]),
    .S(_1119_),
    .Z(_0387_));
 MUX2_X1 _3113_ (.A(pwdata[2]),
    .B(\mem[20] [2]),
    .S(_1119_),
    .Z(_0388_));
 MUX2_X1 _3114_ (.A(pwdata[3]),
    .B(\mem[20] [3]),
    .S(_1119_),
    .Z(_0389_));
 MUX2_X1 _3115_ (.A(pwdata[4]),
    .B(\mem[20] [4]),
    .S(_1119_),
    .Z(_0390_));
 MUX2_X1 _3116_ (.A(pwdata[5]),
    .B(\mem[20] [5]),
    .S(_1119_),
    .Z(_0391_));
 MUX2_X1 _3117_ (.A(pwdata[6]),
    .B(\mem[20] [6]),
    .S(_1119_),
    .Z(_0392_));
 MUX2_X1 _3118_ (.A(pwdata[7]),
    .B(\mem[20] [7]),
    .S(_1119_),
    .Z(_0393_));
 MUX2_X1 _3119_ (.A(pwdata[8]),
    .B(\mem[20] [8]),
    .S(_1119_),
    .Z(_0394_));
 MUX2_X1 _3120_ (.A(pwdata[9]),
    .B(\mem[20] [9]),
    .S(_1119_),
    .Z(_0395_));
 MUX2_X1 _3121_ (.A(pwdata[10]),
    .B(\mem[20] [10]),
    .S(_1119_),
    .Z(_0396_));
 MUX2_X1 _3122_ (.A(pwdata[11]),
    .B(\mem[20] [11]),
    .S(_1119_),
    .Z(_0397_));
 MUX2_X1 _3123_ (.A(pwdata[12]),
    .B(\mem[20] [12]),
    .S(_1119_),
    .Z(_0398_));
 MUX2_X1 _3124_ (.A(pwdata[13]),
    .B(\mem[20] [13]),
    .S(_1119_),
    .Z(_0399_));
 MUX2_X1 _3125_ (.A(pwdata[14]),
    .B(\mem[20] [14]),
    .S(_1119_),
    .Z(_0400_));
 MUX2_X1 _3126_ (.A(pwdata[15]),
    .B(\mem[20] [15]),
    .S(_1119_),
    .Z(_0401_));
 MUX2_X1 _3127_ (.A(pwdata[16]),
    .B(\mem[20] [16]),
    .S(_1119_),
    .Z(_0402_));
 MUX2_X1 _3128_ (.A(pwdata[17]),
    .B(\mem[20] [17]),
    .S(_1119_),
    .Z(_0403_));
 MUX2_X1 _3129_ (.A(pwdata[18]),
    .B(\mem[20] [18]),
    .S(_1119_),
    .Z(_0404_));
 MUX2_X1 _3130_ (.A(pwdata[19]),
    .B(\mem[20] [19]),
    .S(_1119_),
    .Z(_0405_));
 MUX2_X1 _3131_ (.A(pwdata[20]),
    .B(\mem[20] [20]),
    .S(_1119_),
    .Z(_0406_));
 MUX2_X1 _3132_ (.A(pwdata[21]),
    .B(\mem[20] [21]),
    .S(_1119_),
    .Z(_0407_));
 MUX2_X1 _3133_ (.A(pwdata[22]),
    .B(\mem[20] [22]),
    .S(_1119_),
    .Z(_0408_));
 MUX2_X1 _3134_ (.A(pwdata[23]),
    .B(\mem[20] [23]),
    .S(_1119_),
    .Z(_0409_));
 MUX2_X1 _3135_ (.A(pwdata[24]),
    .B(\mem[20] [24]),
    .S(_1119_),
    .Z(_0410_));
 MUX2_X1 _3136_ (.A(pwdata[25]),
    .B(\mem[20] [25]),
    .S(_1119_),
    .Z(_0411_));
 MUX2_X1 _3137_ (.A(pwdata[26]),
    .B(\mem[20] [26]),
    .S(_1119_),
    .Z(_0412_));
 MUX2_X1 _3138_ (.A(pwdata[27]),
    .B(\mem[20] [27]),
    .S(_1119_),
    .Z(_0413_));
 MUX2_X1 _3139_ (.A(pwdata[28]),
    .B(\mem[20] [28]),
    .S(_1119_),
    .Z(_0414_));
 MUX2_X1 _3140_ (.A(pwdata[29]),
    .B(\mem[20] [29]),
    .S(_1119_),
    .Z(_0415_));
 MUX2_X1 _3141_ (.A(pwdata[30]),
    .B(\mem[20] [30]),
    .S(_1119_),
    .Z(_0416_));
 MUX2_X1 _3142_ (.A(pwdata[31]),
    .B(\mem[20] [31]),
    .S(_1119_),
    .Z(_0417_));
 NOR4_X4 _3143_ (.A1(paddr[4]),
    .A2(_1072_),
    .A3(paddr[0]),
    .A4(_1098_),
    .ZN(_1120_));
 NAND2_X4 _3144_ (.A1(_1090_),
    .A2(net50),
    .ZN(_1121_));
 MUX2_X1 _3145_ (.A(pwdata[0]),
    .B(\mem[2] [0]),
    .S(_1121_),
    .Z(_0418_));
 MUX2_X1 _3146_ (.A(pwdata[1]),
    .B(\mem[2] [1]),
    .S(_1121_),
    .Z(_0419_));
 MUX2_X1 _3147_ (.A(pwdata[2]),
    .B(\mem[2] [2]),
    .S(_1121_),
    .Z(_0420_));
 MUX2_X1 _3148_ (.A(pwdata[3]),
    .B(\mem[2] [3]),
    .S(_1121_),
    .Z(_0421_));
 MUX2_X1 _3149_ (.A(pwdata[4]),
    .B(\mem[2] [4]),
    .S(_1121_),
    .Z(_0422_));
 MUX2_X1 _3150_ (.A(pwdata[5]),
    .B(\mem[2] [5]),
    .S(_1121_),
    .Z(_0423_));
 MUX2_X1 _3151_ (.A(pwdata[6]),
    .B(\mem[2] [6]),
    .S(_1121_),
    .Z(_0424_));
 MUX2_X1 _3152_ (.A(pwdata[7]),
    .B(\mem[2] [7]),
    .S(_1121_),
    .Z(_0425_));
 MUX2_X1 _3153_ (.A(pwdata[8]),
    .B(\mem[2] [8]),
    .S(_1121_),
    .Z(_0426_));
 MUX2_X1 _3154_ (.A(pwdata[9]),
    .B(\mem[2] [9]),
    .S(_1121_),
    .Z(_0427_));
 MUX2_X1 _3155_ (.A(pwdata[10]),
    .B(\mem[2] [10]),
    .S(_1121_),
    .Z(_0428_));
 MUX2_X1 _3156_ (.A(pwdata[11]),
    .B(\mem[2] [11]),
    .S(_1121_),
    .Z(_0429_));
 MUX2_X1 _3157_ (.A(pwdata[12]),
    .B(\mem[2] [12]),
    .S(_1121_),
    .Z(_0430_));
 MUX2_X1 _3158_ (.A(pwdata[13]),
    .B(\mem[2] [13]),
    .S(_1121_),
    .Z(_0431_));
 MUX2_X1 _3159_ (.A(pwdata[14]),
    .B(\mem[2] [14]),
    .S(_1121_),
    .Z(_0432_));
 MUX2_X1 _3160_ (.A(pwdata[15]),
    .B(\mem[2] [15]),
    .S(_1121_),
    .Z(_0433_));
 MUX2_X1 _3161_ (.A(pwdata[16]),
    .B(\mem[2] [16]),
    .S(_1121_),
    .Z(_0434_));
 MUX2_X1 _3162_ (.A(pwdata[17]),
    .B(\mem[2] [17]),
    .S(_1121_),
    .Z(_0435_));
 MUX2_X1 _3163_ (.A(pwdata[18]),
    .B(\mem[2] [18]),
    .S(_1121_),
    .Z(_0436_));
 MUX2_X1 _3164_ (.A(pwdata[19]),
    .B(\mem[2] [19]),
    .S(_1121_),
    .Z(_0437_));
 MUX2_X1 _3165_ (.A(pwdata[20]),
    .B(\mem[2] [20]),
    .S(_1121_),
    .Z(_0438_));
 MUX2_X1 _3166_ (.A(pwdata[21]),
    .B(\mem[2] [21]),
    .S(_1121_),
    .Z(_0439_));
 MUX2_X1 _3167_ (.A(pwdata[22]),
    .B(\mem[2] [22]),
    .S(_1121_),
    .Z(_0440_));
 MUX2_X1 _3168_ (.A(pwdata[23]),
    .B(\mem[2] [23]),
    .S(_1121_),
    .Z(_0441_));
 MUX2_X1 _3169_ (.A(pwdata[24]),
    .B(\mem[2] [24]),
    .S(_1121_),
    .Z(_0442_));
 MUX2_X1 _3170_ (.A(pwdata[25]),
    .B(\mem[2] [25]),
    .S(_1121_),
    .Z(_0443_));
 MUX2_X1 _3171_ (.A(pwdata[26]),
    .B(\mem[2] [26]),
    .S(_1121_),
    .Z(_0444_));
 MUX2_X1 _3172_ (.A(pwdata[27]),
    .B(\mem[2] [27]),
    .S(_1121_),
    .Z(_0445_));
 MUX2_X1 _3173_ (.A(pwdata[28]),
    .B(\mem[2] [28]),
    .S(_1121_),
    .Z(_0446_));
 MUX2_X1 _3174_ (.A(pwdata[29]),
    .B(\mem[2] [29]),
    .S(_1121_),
    .Z(_0447_));
 MUX2_X1 _3175_ (.A(pwdata[30]),
    .B(\mem[2] [30]),
    .S(_1121_),
    .Z(_0448_));
 MUX2_X1 _3176_ (.A(pwdata[31]),
    .B(\mem[2] [31]),
    .S(_1121_),
    .Z(_0449_));
 NOR4_X1 _3177_ (.A1(paddr[3]),
    .A2(_1071_),
    .A3(paddr[1]),
    .A4(_1073_),
    .ZN(_1122_));
 AND2_X2 _3178_ (.A1(paddr[4]),
    .A2(_1122_),
    .ZN(_1123_));
 NAND2_X4 _3179_ (.A1(net2),
    .A2(_1123_),
    .ZN(_1124_));
 MUX2_X1 _3180_ (.A(pwdata[0]),
    .B(\mem[21] [0]),
    .S(_1124_),
    .Z(_0450_));
 MUX2_X1 _3181_ (.A(pwdata[1]),
    .B(\mem[21] [1]),
    .S(_1124_),
    .Z(_0451_));
 MUX2_X1 _3182_ (.A(pwdata[2]),
    .B(\mem[21] [2]),
    .S(_1124_),
    .Z(_0452_));
 MUX2_X1 _3183_ (.A(pwdata[3]),
    .B(\mem[21] [3]),
    .S(_1124_),
    .Z(_0453_));
 MUX2_X1 _3184_ (.A(pwdata[4]),
    .B(\mem[21] [4]),
    .S(_1124_),
    .Z(_0454_));
 MUX2_X1 _3185_ (.A(pwdata[5]),
    .B(\mem[21] [5]),
    .S(_1124_),
    .Z(_0455_));
 MUX2_X1 _3186_ (.A(pwdata[6]),
    .B(\mem[21] [6]),
    .S(_1124_),
    .Z(_0456_));
 MUX2_X1 _3187_ (.A(pwdata[7]),
    .B(\mem[21] [7]),
    .S(_1124_),
    .Z(_0457_));
 MUX2_X1 _3188_ (.A(pwdata[8]),
    .B(\mem[21] [8]),
    .S(_1124_),
    .Z(_0458_));
 MUX2_X1 _3189_ (.A(pwdata[9]),
    .B(\mem[21] [9]),
    .S(_1124_),
    .Z(_0459_));
 MUX2_X1 _3190_ (.A(pwdata[10]),
    .B(\mem[21] [10]),
    .S(_1124_),
    .Z(_0460_));
 MUX2_X1 _3191_ (.A(pwdata[11]),
    .B(\mem[21] [11]),
    .S(_1124_),
    .Z(_0461_));
 MUX2_X1 _3192_ (.A(pwdata[12]),
    .B(\mem[21] [12]),
    .S(_1124_),
    .Z(_0462_));
 MUX2_X1 _3193_ (.A(pwdata[13]),
    .B(\mem[21] [13]),
    .S(_1124_),
    .Z(_0463_));
 MUX2_X1 _3194_ (.A(pwdata[14]),
    .B(\mem[21] [14]),
    .S(_1124_),
    .Z(_0464_));
 MUX2_X1 _3195_ (.A(pwdata[15]),
    .B(\mem[21] [15]),
    .S(_1124_),
    .Z(_0465_));
 MUX2_X1 _3196_ (.A(pwdata[16]),
    .B(\mem[21] [16]),
    .S(_1124_),
    .Z(_0466_));
 MUX2_X1 _3197_ (.A(pwdata[17]),
    .B(\mem[21] [17]),
    .S(_1124_),
    .Z(_0467_));
 MUX2_X1 _3198_ (.A(pwdata[18]),
    .B(\mem[21] [18]),
    .S(_1124_),
    .Z(_0468_));
 MUX2_X1 _3199_ (.A(pwdata[19]),
    .B(\mem[21] [19]),
    .S(_1124_),
    .Z(_0469_));
 MUX2_X1 _3200_ (.A(pwdata[20]),
    .B(\mem[21] [20]),
    .S(_1124_),
    .Z(_0470_));
 MUX2_X1 _3201_ (.A(pwdata[21]),
    .B(\mem[21] [21]),
    .S(_1124_),
    .Z(_0471_));
 MUX2_X1 _3202_ (.A(pwdata[22]),
    .B(\mem[21] [22]),
    .S(_1124_),
    .Z(_0472_));
 MUX2_X1 _3203_ (.A(pwdata[23]),
    .B(\mem[21] [23]),
    .S(_1124_),
    .Z(_0473_));
 MUX2_X1 _3204_ (.A(pwdata[24]),
    .B(\mem[21] [24]),
    .S(_1124_),
    .Z(_0474_));
 MUX2_X1 _3205_ (.A(pwdata[25]),
    .B(\mem[21] [25]),
    .S(_1124_),
    .Z(_0475_));
 MUX2_X1 _3206_ (.A(pwdata[26]),
    .B(\mem[21] [26]),
    .S(_1124_),
    .Z(_0476_));
 MUX2_X1 _3207_ (.A(pwdata[27]),
    .B(\mem[21] [27]),
    .S(_1124_),
    .Z(_0477_));
 MUX2_X1 _3208_ (.A(pwdata[28]),
    .B(\mem[21] [28]),
    .S(_1124_),
    .Z(_0478_));
 MUX2_X1 _3209_ (.A(pwdata[29]),
    .B(\mem[21] [29]),
    .S(_1124_),
    .Z(_0479_));
 MUX2_X1 _3210_ (.A(pwdata[30]),
    .B(\mem[21] [30]),
    .S(_1124_),
    .Z(_0480_));
 MUX2_X1 _3211_ (.A(pwdata[31]),
    .B(\mem[21] [31]),
    .S(_1124_),
    .Z(_0481_));
 NOR4_X4 _3212_ (.A1(_1069_),
    .A2(_1072_),
    .A3(paddr[0]),
    .A4(_1075_),
    .ZN(_1125_));
 NAND2_X4 _3213_ (.A1(net2),
    .A2(net48),
    .ZN(_1126_));
 MUX2_X1 _3214_ (.A(pwdata[0]),
    .B(\mem[30] [0]),
    .S(_1126_),
    .Z(_0482_));
 MUX2_X1 _3215_ (.A(pwdata[1]),
    .B(\mem[30] [1]),
    .S(_1126_),
    .Z(_0483_));
 MUX2_X1 _3216_ (.A(pwdata[2]),
    .B(\mem[30] [2]),
    .S(_1126_),
    .Z(_0484_));
 MUX2_X1 _3217_ (.A(pwdata[3]),
    .B(\mem[30] [3]),
    .S(_1126_),
    .Z(_0485_));
 MUX2_X1 _3218_ (.A(pwdata[4]),
    .B(\mem[30] [4]),
    .S(_1126_),
    .Z(_0486_));
 MUX2_X1 _3219_ (.A(pwdata[5]),
    .B(\mem[30] [5]),
    .S(_1126_),
    .Z(_0487_));
 MUX2_X1 _3220_ (.A(pwdata[6]),
    .B(\mem[30] [6]),
    .S(_1126_),
    .Z(_0488_));
 MUX2_X1 _3221_ (.A(pwdata[7]),
    .B(\mem[30] [7]),
    .S(_1126_),
    .Z(_0489_));
 MUX2_X1 _3222_ (.A(pwdata[8]),
    .B(\mem[30] [8]),
    .S(_1126_),
    .Z(_0490_));
 MUX2_X1 _3223_ (.A(pwdata[9]),
    .B(\mem[30] [9]),
    .S(_1126_),
    .Z(_0491_));
 MUX2_X1 _3224_ (.A(pwdata[10]),
    .B(\mem[30] [10]),
    .S(_1126_),
    .Z(_0492_));
 MUX2_X1 _3225_ (.A(pwdata[11]),
    .B(\mem[30] [11]),
    .S(_1126_),
    .Z(_0493_));
 MUX2_X1 _3226_ (.A(pwdata[12]),
    .B(\mem[30] [12]),
    .S(_1126_),
    .Z(_0494_));
 MUX2_X1 _3227_ (.A(pwdata[13]),
    .B(\mem[30] [13]),
    .S(_1126_),
    .Z(_0495_));
 MUX2_X1 _3228_ (.A(pwdata[14]),
    .B(\mem[30] [14]),
    .S(_1126_),
    .Z(_0496_));
 MUX2_X1 _3229_ (.A(pwdata[15]),
    .B(\mem[30] [15]),
    .S(_1126_),
    .Z(_0497_));
 MUX2_X1 _3230_ (.A(pwdata[16]),
    .B(\mem[30] [16]),
    .S(_1126_),
    .Z(_0498_));
 MUX2_X1 _3231_ (.A(pwdata[17]),
    .B(\mem[30] [17]),
    .S(_1126_),
    .Z(_0499_));
 MUX2_X1 _3232_ (.A(pwdata[18]),
    .B(\mem[30] [18]),
    .S(_1126_),
    .Z(_0500_));
 MUX2_X1 _3233_ (.A(pwdata[19]),
    .B(\mem[30] [19]),
    .S(_1126_),
    .Z(_0501_));
 MUX2_X1 _3234_ (.A(pwdata[20]),
    .B(\mem[30] [20]),
    .S(_1126_),
    .Z(_0502_));
 MUX2_X1 _3235_ (.A(pwdata[21]),
    .B(\mem[30] [21]),
    .S(_1126_),
    .Z(_0503_));
 MUX2_X1 _3236_ (.A(pwdata[22]),
    .B(\mem[30] [22]),
    .S(_1126_),
    .Z(_0504_));
 MUX2_X1 _3237_ (.A(pwdata[23]),
    .B(\mem[30] [23]),
    .S(_1126_),
    .Z(_0505_));
 MUX2_X1 _3238_ (.A(pwdata[24]),
    .B(\mem[30] [24]),
    .S(_1126_),
    .Z(_0506_));
 MUX2_X1 _3239_ (.A(pwdata[25]),
    .B(\mem[30] [25]),
    .S(_1126_),
    .Z(_0507_));
 MUX2_X1 _3240_ (.A(pwdata[26]),
    .B(\mem[30] [26]),
    .S(_1126_),
    .Z(_0508_));
 MUX2_X1 _3241_ (.A(pwdata[27]),
    .B(\mem[30] [27]),
    .S(_1126_),
    .Z(_0509_));
 MUX2_X1 _3242_ (.A(pwdata[28]),
    .B(\mem[30] [28]),
    .S(_1126_),
    .Z(_0510_));
 MUX2_X1 _3243_ (.A(pwdata[29]),
    .B(\mem[30] [29]),
    .S(_1126_),
    .Z(_0511_));
 MUX2_X1 _3244_ (.A(pwdata[30]),
    .B(\mem[30] [30]),
    .S(_1126_),
    .Z(_0512_));
 MUX2_X1 _3245_ (.A(pwdata[31]),
    .B(\mem[30] [31]),
    .S(_1126_),
    .Z(_0513_));
 NOR4_X1 _3246_ (.A1(paddr[3]),
    .A2(_1071_),
    .A3(_1072_),
    .A4(paddr[0]),
    .ZN(_1127_));
 AND2_X2 _3247_ (.A1(paddr[4]),
    .A2(_1127_),
    .ZN(_1128_));
 NAND2_X4 _3248_ (.A1(_1090_),
    .A2(_1128_),
    .ZN(_1129_));
 MUX2_X1 _3249_ (.A(pwdata[0]),
    .B(\mem[22] [0]),
    .S(_1129_),
    .Z(_0514_));
 MUX2_X1 _3250_ (.A(pwdata[1]),
    .B(\mem[22] [1]),
    .S(_1129_),
    .Z(_0515_));
 MUX2_X1 _3251_ (.A(pwdata[2]),
    .B(\mem[22] [2]),
    .S(_1129_),
    .Z(_0516_));
 MUX2_X1 _3252_ (.A(pwdata[3]),
    .B(\mem[22] [3]),
    .S(_1129_),
    .Z(_0517_));
 MUX2_X1 _3253_ (.A(pwdata[4]),
    .B(\mem[22] [4]),
    .S(_1129_),
    .Z(_0518_));
 MUX2_X1 _3254_ (.A(pwdata[5]),
    .B(\mem[22] [5]),
    .S(_1129_),
    .Z(_0519_));
 MUX2_X1 _3255_ (.A(pwdata[6]),
    .B(\mem[22] [6]),
    .S(_1129_),
    .Z(_0520_));
 MUX2_X1 _3256_ (.A(pwdata[7]),
    .B(\mem[22] [7]),
    .S(_1129_),
    .Z(_0521_));
 MUX2_X1 _3257_ (.A(pwdata[8]),
    .B(\mem[22] [8]),
    .S(_1129_),
    .Z(_0522_));
 MUX2_X1 _3258_ (.A(pwdata[9]),
    .B(\mem[22] [9]),
    .S(_1129_),
    .Z(_0523_));
 MUX2_X1 _3259_ (.A(pwdata[10]),
    .B(\mem[22] [10]),
    .S(_1129_),
    .Z(_0524_));
 MUX2_X1 _3260_ (.A(pwdata[11]),
    .B(\mem[22] [11]),
    .S(_1129_),
    .Z(_0525_));
 MUX2_X1 _3261_ (.A(pwdata[12]),
    .B(\mem[22] [12]),
    .S(_1129_),
    .Z(_0526_));
 MUX2_X1 _3262_ (.A(pwdata[13]),
    .B(\mem[22] [13]),
    .S(_1129_),
    .Z(_0527_));
 MUX2_X1 _3263_ (.A(pwdata[14]),
    .B(\mem[22] [14]),
    .S(_1129_),
    .Z(_0528_));
 MUX2_X1 _3264_ (.A(pwdata[15]),
    .B(\mem[22] [15]),
    .S(_1129_),
    .Z(_0529_));
 MUX2_X1 _3265_ (.A(pwdata[16]),
    .B(\mem[22] [16]),
    .S(_1129_),
    .Z(_0530_));
 MUX2_X1 _3266_ (.A(pwdata[17]),
    .B(\mem[22] [17]),
    .S(_1129_),
    .Z(_0531_));
 MUX2_X1 _3267_ (.A(pwdata[18]),
    .B(\mem[22] [18]),
    .S(_1129_),
    .Z(_0532_));
 MUX2_X1 _3268_ (.A(pwdata[19]),
    .B(\mem[22] [19]),
    .S(_1129_),
    .Z(_0533_));
 MUX2_X1 _3269_ (.A(pwdata[20]),
    .B(\mem[22] [20]),
    .S(_1129_),
    .Z(_0534_));
 MUX2_X1 _3270_ (.A(pwdata[21]),
    .B(\mem[22] [21]),
    .S(_1129_),
    .Z(_0535_));
 MUX2_X1 _3271_ (.A(pwdata[22]),
    .B(\mem[22] [22]),
    .S(_1129_),
    .Z(_0536_));
 MUX2_X1 _3272_ (.A(pwdata[23]),
    .B(\mem[22] [23]),
    .S(_1129_),
    .Z(_0537_));
 MUX2_X1 _3273_ (.A(pwdata[24]),
    .B(\mem[22] [24]),
    .S(_1129_),
    .Z(_0538_));
 MUX2_X1 _3274_ (.A(pwdata[25]),
    .B(\mem[22] [25]),
    .S(_1129_),
    .Z(_0539_));
 MUX2_X1 _3275_ (.A(pwdata[26]),
    .B(\mem[22] [26]),
    .S(_1129_),
    .Z(_0540_));
 MUX2_X1 _3276_ (.A(pwdata[27]),
    .B(\mem[22] [27]),
    .S(_1129_),
    .Z(_0541_));
 MUX2_X1 _3277_ (.A(pwdata[28]),
    .B(\mem[22] [28]),
    .S(_1129_),
    .Z(_0542_));
 MUX2_X1 _3278_ (.A(pwdata[29]),
    .B(\mem[22] [29]),
    .S(_1129_),
    .Z(_0543_));
 MUX2_X1 _3279_ (.A(pwdata[30]),
    .B(\mem[22] [30]),
    .S(_1129_),
    .Z(_0544_));
 MUX2_X1 _3280_ (.A(pwdata[31]),
    .B(\mem[22] [31]),
    .S(_1129_),
    .Z(_0545_));
 AND3_X2 _3281_ (.A1(_1074_),
    .A2(penable),
    .A3(_2855_[0]),
    .ZN(_1130_));
 NAND3_X2 _3282_ (.A1(_1074_),
    .A2(penable),
    .A3(_2855_[0]),
    .ZN(_1131_));
 NOR2_X1 _3283_ (.A1(prdata[0]),
    .A2(_1130_),
    .ZN(_1132_));
 NOR3_X4 _3284_ (.A1(paddr[4]),
    .A2(_1076_),
    .A3(_1098_),
    .ZN(_1133_));
 NOR3_X4 _3285_ (.A1(paddr[4]),
    .A2(_1092_),
    .A3(_1098_),
    .ZN(_1134_));
 AND2_X2 _3286_ (.A1(_1069_),
    .A2(_1095_),
    .ZN(_1135_));
 AOI22_X1 _3287_ (.A1(\mem[20] [0]),
    .A2(net53),
    .B1(net51),
    .B2(\mem[2] [0]),
    .ZN(_1136_));
 NOR4_X4 _3288_ (.A1(paddr[4]),
    .A2(paddr[3]),
    .A3(_1071_),
    .A4(_1076_),
    .ZN(_1137_));
 AND2_X2 _3289_ (.A1(_1069_),
    .A2(_1122_),
    .ZN(_1138_));
 NOR4_X4 _3290_ (.A1(paddr[4]),
    .A2(_1070_),
    .A3(paddr[2]),
    .A4(_1092_),
    .ZN(_1139_));
 NOR4_X4 _3291_ (.A1(_1069_),
    .A2(paddr[3]),
    .A3(_1071_),
    .A4(_1092_),
    .ZN(_1140_));
 NOR4_X4 _3292_ (.A1(paddr[4]),
    .A2(paddr[1]),
    .A3(_1073_),
    .A4(_1075_),
    .ZN(_1141_));
 NOR4_X4 _3293_ (.A1(paddr[4]),
    .A2(_1072_),
    .A3(paddr[0]),
    .A4(_1075_),
    .ZN(_1142_));
 NOR4_X4 _3294_ (.A1(_1069_),
    .A2(paddr[1]),
    .A3(_1073_),
    .A4(_1075_),
    .ZN(_1143_));
 AOI22_X1 _3295_ (.A1(\mem[18] [0]),
    .A2(net63),
    .B1(net59),
    .B2(\mem[19] [0]),
    .ZN(_1144_));
 NOR4_X4 _3296_ (.A1(paddr[4]),
    .A2(paddr[1]),
    .A3(_1073_),
    .A4(_1098_),
    .ZN(_1145_));
 AND2_X2 _3297_ (.A1(paddr[4]),
    .A2(_1115_),
    .ZN(_1146_));
 AND2_X2 _3298_ (.A1(_1069_),
    .A2(_1127_),
    .ZN(_1147_));
 NOR4_X4 _3299_ (.A1(paddr[4]),
    .A2(_1070_),
    .A3(paddr[2]),
    .A4(_1076_),
    .ZN(_1148_));
 NOR4_X4 _3300_ (.A1(paddr[4]),
    .A2(paddr[3]),
    .A3(_1071_),
    .A4(_1092_),
    .ZN(_1149_));
 AOI222_X2 _3301_ (.A1(\mem[15] [0]),
    .A2(net12),
    .B1(_1128_),
    .B2(\mem[22] [0]),
    .C1(net31),
    .C2(\mem[13] [0]),
    .ZN(_1150_));
 AOI221_X1 _3302_ (.A(_1131_),
    .B1(net37),
    .B2(\mem[11] [0]),
    .C1(net35),
    .C2(\mem[23] [0]),
    .ZN(_1151_));
 NAND2_X1 _3303_ (.A1(_1150_),
    .A2(_1151_),
    .ZN(_1152_));
 AOI22_X1 _3304_ (.A1(\mem[17] [0]),
    .A2(net70),
    .B1(_1123_),
    .B2(\mem[21] [0]),
    .ZN(_1153_));
 AOI22_X1 _3305_ (.A1(\mem[14] [0]),
    .A2(net28),
    .B1(net20),
    .B2(\mem[8] [0]),
    .ZN(_1154_));
 AOI22_X1 _3306_ (.A1(\mem[5] [0]),
    .A2(_1138_),
    .B1(_1146_),
    .B2(\mem[25] [0]),
    .ZN(_1155_));
 NAND4_X1 _3307_ (.A1(_1136_),
    .A2(_1153_),
    .A3(_1154_),
    .A4(_1155_),
    .ZN(_1156_));
 NOR2_X1 _3308_ (.A1(_1152_),
    .A2(_1156_),
    .ZN(_1157_));
 AOI222_X1 _3309_ (.A1(\mem[4] [0]),
    .A2(net41),
    .B1(_1147_),
    .B2(\mem[6] [0]),
    .C1(net23),
    .C2(\mem[1] [0]),
    .ZN(_1158_));
 AOI222_X1 _3310_ (.A1(\mem[28] [0]),
    .A2(net62),
    .B1(net56),
    .B2(\mem[24] [0]),
    .C1(net16),
    .C2(\mem[7] [0]),
    .ZN(_1159_));
 AOI222_X1 _3311_ (.A1(\mem[31] [0]),
    .A2(net7),
    .B1(net48),
    .B2(\mem[30] [0]),
    .C1(net26),
    .C2(\mem[29] [0]),
    .ZN(_1160_));
 NAND4_X1 _3312_ (.A1(_1144_),
    .A2(_1158_),
    .A3(_1159_),
    .A4(_1160_),
    .ZN(_1161_));
 AOI22_X1 _3313_ (.A1(\mem[0] [0]),
    .A2(net45),
    .B1(net43),
    .B2(\mem[3] [0]),
    .ZN(_1162_));
 AOI22_X1 _3314_ (.A1(\mem[12] [0]),
    .A2(net15),
    .B1(net9),
    .B2(\mem[16] [0]),
    .ZN(_1163_));
 AOI22_X1 _3315_ (.A1(\mem[9] [0]),
    .A2(net5),
    .B1(_1135_),
    .B2(\mem[10] [0]),
    .ZN(_1164_));
 AOI22_X1 _3316_ (.A1(\mem[26] [0]),
    .A2(_1096_),
    .B1(_1105_),
    .B2(\mem[27] [0]),
    .ZN(_1165_));
 NAND4_X1 _3317_ (.A1(_1162_),
    .A2(_1163_),
    .A3(_1164_),
    .A4(_1165_),
    .ZN(_1166_));
 NOR2_X1 _3318_ (.A1(_1161_),
    .A2(_1166_),
    .ZN(_1167_));
 AOI21_X1 _3319_ (.A(_1132_),
    .B1(_1157_),
    .B2(_1167_),
    .ZN(_0546_));
 AOI22_X1 _3320_ (.A1(\mem[18] [1]),
    .A2(net64),
    .B1(net60),
    .B2(\mem[19] [1]),
    .ZN(_1168_));
 AOI222_X1 _3321_ (.A1(\mem[16] [1]),
    .A2(net11),
    .B1(_1123_),
    .B2(\mem[21] [1]),
    .C1(_1146_),
    .C2(\mem[25] [1]),
    .ZN(_1169_));
 AOI221_X1 _3322_ (.A(net4),
    .B1(net55),
    .B2(\mem[20] [1]),
    .C1(\mem[12] [1]),
    .C2(net15),
    .ZN(_1170_));
 AOI22_X1 _3323_ (.A1(\mem[15] [1]),
    .A2(net12),
    .B1(net61),
    .B2(\mem[28] [1]),
    .ZN(_1171_));
 AOI22_X1 _3324_ (.A1(\mem[17] [1]),
    .A2(net68),
    .B1(_1143_),
    .B2(\mem[29] [1]),
    .ZN(_1172_));
 AOI22_X1 _3325_ (.A1(\mem[4] [1]),
    .A2(net40),
    .B1(net17),
    .B2(\mem[7] [1]),
    .ZN(_1173_));
 AND4_X1 _3326_ (.A1(_1168_),
    .A2(_1171_),
    .A3(_1172_),
    .A4(_1173_),
    .ZN(_1174_));
 NAND3_X1 _3327_ (.A1(_1169_),
    .A2(_1170_),
    .A3(_1174_),
    .ZN(_1175_));
 AOI22_X1 _3328_ (.A1(\mem[26] [1]),
    .A2(_1096_),
    .B1(net66),
    .B2(\mem[27] [1]),
    .ZN(_1176_));
 AOI222_X1 _3329_ (.A1(\mem[0] [1]),
    .A2(net45),
    .B1(_1138_),
    .B2(\mem[5] [1]),
    .C1(\mem[1] [1]),
    .C2(net24),
    .ZN(_1177_));
 AOI222_X1 _3330_ (.A1(\mem[9] [1]),
    .A2(net6),
    .B1(_1135_),
    .B2(\mem[10] [1]),
    .C1(_1147_),
    .C2(\mem[6] [1]),
    .ZN(_1178_));
 AOI222_X1 _3331_ (.A1(\mem[31] [1]),
    .A2(_1101_),
    .B1(net56),
    .B2(\mem[24] [1]),
    .C1(net47),
    .C2(\mem[30] [1]),
    .ZN(_1179_));
 NAND4_X1 _3332_ (.A1(_1176_),
    .A2(_1177_),
    .A3(_1178_),
    .A4(_1179_),
    .ZN(_1180_));
 AOI22_X1 _3333_ (.A1(\mem[14] [1]),
    .A2(net27),
    .B1(net21),
    .B2(\mem[8] [1]),
    .ZN(_1181_));
 AOI22_X1 _3334_ (.A1(\mem[22] [1]),
    .A2(_1128_),
    .B1(net37),
    .B2(\mem[11] [1]),
    .ZN(_1182_));
 AOI22_X1 _3335_ (.A1(\mem[2] [1]),
    .A2(net51),
    .B1(net36),
    .B2(\mem[23] [1]),
    .ZN(_1183_));
 AOI22_X1 _3336_ (.A1(\mem[3] [1]),
    .A2(net44),
    .B1(net32),
    .B2(\mem[13] [1]),
    .ZN(_1184_));
 NAND4_X1 _3337_ (.A1(_1181_),
    .A2(_1182_),
    .A3(_1183_),
    .A4(_1184_),
    .ZN(_1185_));
 NOR3_X1 _3338_ (.A1(_1175_),
    .A2(_1180_),
    .A3(_1185_),
    .ZN(_1186_));
 AOI21_X1 _3339_ (.A(_1186_),
    .B1(net4),
    .B2(_1059_),
    .ZN(_0547_));
 AOI22_X1 _3340_ (.A1(\mem[22] [2]),
    .A2(_1128_),
    .B1(net37),
    .B2(\mem[11] [2]),
    .ZN(_1187_));
 AOI22_X1 _3341_ (.A1(\mem[14] [2]),
    .A2(net29),
    .B1(net20),
    .B2(\mem[8] [2]),
    .ZN(_1188_));
 AOI22_X1 _3342_ (.A1(\mem[4] [2]),
    .A2(net42),
    .B1(net36),
    .B2(\mem[23] [2]),
    .ZN(_1189_));
 AOI22_X1 _3343_ (.A1(\mem[12] [2]),
    .A2(_1077_),
    .B1(net43),
    .B2(\mem[3] [2]),
    .ZN(_1190_));
 NAND4_X1 _3344_ (.A1(_1187_),
    .A2(_1188_),
    .A3(_1189_),
    .A4(_1190_),
    .ZN(_1191_));
 AOI22_X1 _3345_ (.A1(\mem[26] [2]),
    .A2(_1096_),
    .B1(_1105_),
    .B2(\mem[27] [2]),
    .ZN(_1192_));
 AOI222_X1 _3346_ (.A1(\mem[5] [2]),
    .A2(_1138_),
    .B1(_1147_),
    .B2(\mem[6] [2]),
    .C1(net23),
    .C2(\mem[1] [2]),
    .ZN(_1193_));
 AOI222_X1 _3347_ (.A1(\mem[9] [2]),
    .A2(net5),
    .B1(_1135_),
    .B2(\mem[10] [2]),
    .C1(net18),
    .C2(\mem[7] [2]),
    .ZN(_1194_));
 AOI222_X1 _3348_ (.A1(\mem[31] [2]),
    .A2(net7),
    .B1(net57),
    .B2(\mem[24] [2]),
    .C1(net49),
    .C2(\mem[30] [2]),
    .ZN(_1195_));
 NAND4_X1 _3349_ (.A1(_1192_),
    .A2(_1193_),
    .A3(_1194_),
    .A4(_1195_),
    .ZN(_1196_));
 AOI222_X1 _3350_ (.A1(\mem[16] [2]),
    .A2(net9),
    .B1(_1123_),
    .B2(\mem[21] [2]),
    .C1(_1146_),
    .C2(\mem[25] [2]),
    .ZN(_1197_));
 AOI221_X1 _3351_ (.A(net3),
    .B1(net34),
    .B2(\mem[13] [2]),
    .C1(net53),
    .C2(\mem[20] [2]),
    .ZN(_1198_));
 AOI22_X1 _3352_ (.A1(\mem[18] [2]),
    .A2(net63),
    .B1(net60),
    .B2(\mem[19] [2]),
    .ZN(_1199_));
 AOI22_X1 _3353_ (.A1(\mem[15] [2]),
    .A2(net12),
    .B1(net61),
    .B2(\mem[28] [2]),
    .ZN(_1200_));
 AOI22_X1 _3354_ (.A1(\mem[17] [2]),
    .A2(net68),
    .B1(net26),
    .B2(\mem[29] [2]),
    .ZN(_1201_));
 AOI22_X1 _3355_ (.A1(\mem[2] [2]),
    .A2(net51),
    .B1(net45),
    .B2(\mem[0] [2]),
    .ZN(_1202_));
 AND4_X1 _3356_ (.A1(_1199_),
    .A2(_1200_),
    .A3(_1201_),
    .A4(_1202_),
    .ZN(_1203_));
 NAND3_X1 _3357_ (.A1(_1197_),
    .A2(_1198_),
    .A3(_1203_),
    .ZN(_1204_));
 NOR3_X1 _3358_ (.A1(_1191_),
    .A2(_1196_),
    .A3(_1204_),
    .ZN(_1205_));
 AOI21_X1 _3359_ (.A(_1205_),
    .B1(net3),
    .B2(_1060_),
    .ZN(_0548_));
 NOR2_X1 _3360_ (.A1(prdata[3]),
    .A2(_1130_),
    .ZN(_1206_));
 AOI22_X1 _3361_ (.A1(\mem[2] [3]),
    .A2(net50),
    .B1(_1134_),
    .B2(\mem[3] [3]),
    .ZN(_1207_));
 AOI222_X1 _3362_ (.A1(\mem[17] [3]),
    .A2(net69),
    .B1(_1123_),
    .B2(\mem[21] [3]),
    .C1(_1128_),
    .C2(\mem[22] [3]),
    .ZN(_1208_));
 AOI221_X1 _3363_ (.A(_1131_),
    .B1(_1147_),
    .B2(\mem[6] [3]),
    .C1(net10),
    .C2(\mem[16] [3]),
    .ZN(_1209_));
 NAND2_X1 _3364_ (.A1(_1208_),
    .A2(_1209_),
    .ZN(_1210_));
 AOI22_X1 _3365_ (.A1(\mem[27] [3]),
    .A2(net67),
    .B1(net16),
    .B2(\mem[7] [3]),
    .ZN(_1211_));
 AOI22_X1 _3366_ (.A1(\mem[26] [3]),
    .A2(_1096_),
    .B1(_1146_),
    .B2(\mem[25] [3]),
    .ZN(_1212_));
 AOI22_X1 _3367_ (.A1(\mem[15] [3]),
    .A2(net13),
    .B1(net33),
    .B2(\mem[13] [3]),
    .ZN(_1213_));
 NAND4_X1 _3368_ (.A1(_1207_),
    .A2(_1211_),
    .A3(_1212_),
    .A4(_1213_),
    .ZN(_1214_));
 NOR2_X1 _3369_ (.A1(_1210_),
    .A2(_1214_),
    .ZN(_1215_));
 AOI22_X1 _3370_ (.A1(\mem[18] [3]),
    .A2(net65),
    .B1(net59),
    .B2(\mem[19] [3]),
    .ZN(_1216_));
 AOI222_X2 _3371_ (.A1(\mem[12] [3]),
    .A2(net14),
    .B1(net29),
    .B2(\mem[14] [3]),
    .C1(net19),
    .C2(\mem[8] [3]),
    .ZN(_1217_));
 AOI222_X1 _3372_ (.A1(\mem[28] [3]),
    .A2(net62),
    .B1(net58),
    .B2(\mem[24] [3]),
    .C1(net5),
    .C2(\mem[9] [3]),
    .ZN(_1218_));
 AOI222_X1 _3373_ (.A1(\mem[31] [3]),
    .A2(net8),
    .B1(net48),
    .B2(\mem[30] [3]),
    .C1(net25),
    .C2(\mem[29] [3]),
    .ZN(_1219_));
 NAND4_X1 _3374_ (.A1(_1216_),
    .A2(_1217_),
    .A3(_1218_),
    .A4(_1219_),
    .ZN(_1220_));
 AOI22_X1 _3375_ (.A1(\mem[4] [3]),
    .A2(net42),
    .B1(net23),
    .B2(\mem[1] [3]),
    .ZN(_1221_));
 AOI22_X1 _3376_ (.A1(\mem[20] [3]),
    .A2(net54),
    .B1(net46),
    .B2(\mem[0] [3]),
    .ZN(_1222_));
 AOI22_X1 _3377_ (.A1(\mem[10] [3]),
    .A2(_1135_),
    .B1(_1138_),
    .B2(\mem[5] [3]),
    .ZN(_1223_));
 AOI22_X1 _3378_ (.A1(\mem[11] [3]),
    .A2(net38),
    .B1(net35),
    .B2(\mem[23] [3]),
    .ZN(_1224_));
 NAND4_X1 _3379_ (.A1(_1221_),
    .A2(_1222_),
    .A3(_1223_),
    .A4(_1224_),
    .ZN(_1225_));
 NOR2_X1 _3380_ (.A1(_1220_),
    .A2(_1225_),
    .ZN(_1226_));
 AOI21_X1 _3381_ (.A(_1206_),
    .B1(_1215_),
    .B2(_1226_),
    .ZN(_0549_));
 AOI222_X1 _3382_ (.A1(\mem[4] [4]),
    .A2(net41),
    .B1(_1147_),
    .B2(\mem[6] [4]),
    .C1(net24),
    .C2(\mem[1] [4]),
    .ZN(_1227_));
 AOI22_X1 _3383_ (.A1(\mem[26] [4]),
    .A2(_1096_),
    .B1(net44),
    .B2(\mem[3] [4]),
    .ZN(_1228_));
 AOI222_X1 _3384_ (.A1(\mem[15] [4]),
    .A2(net12),
    .B1(net53),
    .B2(\mem[20] [4]),
    .C1(_1128_),
    .C2(\mem[22] [4]),
    .ZN(_1229_));
 AOI222_X1 _3385_ (.A1(\mem[16] [4]),
    .A2(net9),
    .B1(_1105_),
    .B2(\mem[27] [4]),
    .C1(net51),
    .C2(\mem[2] [4]),
    .ZN(_1230_));
 NAND4_X1 _3386_ (.A1(_1227_),
    .A2(_1228_),
    .A3(_1229_),
    .A4(_1230_),
    .ZN(_1231_));
 AOI22_X1 _3387_ (.A1(\mem[28] [4]),
    .A2(net61),
    .B1(_1138_),
    .B2(\mem[5] [4]),
    .ZN(_1232_));
 AOI222_X1 _3388_ (.A1(\mem[31] [4]),
    .A2(net7),
    .B1(net45),
    .B2(\mem[0] [4]),
    .C1(net18),
    .C2(\mem[7] [4]),
    .ZN(_1233_));
 AOI221_X1 _3389_ (.A(net4),
    .B1(net37),
    .B2(\mem[11] [4]),
    .C1(net21),
    .C2(\mem[8] [4]),
    .ZN(_1234_));
 AOI222_X2 _3390_ (.A1(\mem[24] [4]),
    .A2(net56),
    .B1(_1135_),
    .B2(\mem[10] [4]),
    .C1(net31),
    .C2(\mem[13] [4]),
    .ZN(_1235_));
 NAND4_X1 _3391_ (.A1(_1232_),
    .A2(_1233_),
    .A3(_1234_),
    .A4(_1235_),
    .ZN(_1236_));
 AOI22_X1 _3392_ (.A1(\mem[18] [4]),
    .A2(net63),
    .B1(net60),
    .B2(\mem[19] [4]),
    .ZN(_1237_));
 AOI222_X1 _3393_ (.A1(\mem[17] [4]),
    .A2(net70),
    .B1(_1123_),
    .B2(\mem[21] [4]),
    .C1(net36),
    .C2(\mem[23] [4]),
    .ZN(_1238_));
 AOI222_X2 _3394_ (.A1(\mem[12] [4]),
    .A2(net15),
    .B1(net5),
    .B2(\mem[9] [4]),
    .C1(net28),
    .C2(\mem[14] [4]),
    .ZN(_1239_));
 NAND3_X1 _3395_ (.A1(_1237_),
    .A2(_1238_),
    .A3(_1239_),
    .ZN(_1240_));
 AOI222_X1 _3396_ (.A1(\mem[30] [4]),
    .A2(net47),
    .B1(net26),
    .B2(\mem[29] [4]),
    .C1(_1146_),
    .C2(\mem[25] [4]),
    .ZN(_1241_));
 INV_X1 _3397_ (.A(_1241_),
    .ZN(_1242_));
 NOR4_X1 _3398_ (.A1(_1231_),
    .A2(_1236_),
    .A3(_1240_),
    .A4(_1242_),
    .ZN(_1243_));
 AOI21_X1 _3399_ (.A(_1243_),
    .B1(net4),
    .B2(_1061_),
    .ZN(_0550_));
 NOR2_X1 _3400_ (.A1(prdata[5]),
    .A2(_1130_),
    .ZN(_1244_));
 AOI22_X1 _3401_ (.A1(\mem[0] [5]),
    .A2(net46),
    .B1(net35),
    .B2(\mem[23] [5]),
    .ZN(_1245_));
 AOI22_X1 _3402_ (.A1(\mem[4] [5]),
    .A2(net42),
    .B1(net23),
    .B2(\mem[1] [5]),
    .ZN(_1246_));
 AOI22_X1 _3403_ (.A1(\mem[10] [5]),
    .A2(_1135_),
    .B1(_1138_),
    .B2(\mem[5] [5]),
    .ZN(_1247_));
 AOI22_X1 _3404_ (.A1(\mem[20] [5]),
    .A2(net54),
    .B1(net38),
    .B2(\mem[11] [5]),
    .ZN(_1248_));
 AND4_X1 _3405_ (.A1(_1245_),
    .A2(_1246_),
    .A3(_1247_),
    .A4(_1248_),
    .ZN(_1249_));
 AOI22_X1 _3406_ (.A1(\mem[18] [5]),
    .A2(net65),
    .B1(net60),
    .B2(\mem[19] [5]),
    .ZN(_1250_));
 AOI222_X2 _3407_ (.A1(\mem[9] [5]),
    .A2(net5),
    .B1(net33),
    .B2(\mem[13] [5]),
    .C1(net22),
    .C2(\mem[8] [5]),
    .ZN(_1251_));
 AOI222_X2 _3408_ (.A1(\mem[28] [5]),
    .A2(_1109_),
    .B1(net58),
    .B2(\mem[24] [5]),
    .C1(net30),
    .C2(\mem[14] [5]),
    .ZN(_1252_));
 AOI222_X1 _3409_ (.A1(\mem[31] [5]),
    .A2(net8),
    .B1(net49),
    .B2(\mem[30] [5]),
    .C1(net25),
    .C2(\mem[29] [5]),
    .ZN(_1253_));
 NAND4_X1 _3410_ (.A1(_1250_),
    .A2(_1251_),
    .A3(_1252_),
    .A4(_1253_),
    .ZN(_1254_));
 AOI222_X1 _3411_ (.A1(\mem[17] [5]),
    .A2(net69),
    .B1(_1123_),
    .B2(\mem[21] [5]),
    .C1(_1128_),
    .C2(\mem[22] [5]),
    .ZN(_1255_));
 AOI221_X1 _3412_ (.A(_1131_),
    .B1(_1147_),
    .B2(\mem[6] [5]),
    .C1(net10),
    .C2(\mem[16] [5]),
    .ZN(_1256_));
 NAND2_X1 _3413_ (.A1(_1255_),
    .A2(_1256_),
    .ZN(_1257_));
 AOI22_X1 _3414_ (.A1(\mem[2] [5]),
    .A2(net50),
    .B1(_1134_),
    .B2(\mem[3] [5]),
    .ZN(_1258_));
 AOI22_X1 _3415_ (.A1(\mem[27] [5]),
    .A2(net67),
    .B1(net16),
    .B2(\mem[7] [5]),
    .ZN(_1259_));
 AOI22_X1 _3416_ (.A1(\mem[26] [5]),
    .A2(_1096_),
    .B1(_1146_),
    .B2(\mem[25] [5]),
    .ZN(_1260_));
 AOI22_X1 _3417_ (.A1(\mem[12] [5]),
    .A2(net14),
    .B1(net13),
    .B2(\mem[15] [5]),
    .ZN(_1261_));
 NAND4_X1 _3418_ (.A1(_1258_),
    .A2(_1259_),
    .A3(_1260_),
    .A4(_1261_),
    .ZN(_1262_));
 NOR3_X1 _3419_ (.A1(_1254_),
    .A2(_1257_),
    .A3(_1262_),
    .ZN(_1263_));
 AOI21_X1 _3420_ (.A(_1244_),
    .B1(_1249_),
    .B2(_1263_),
    .ZN(_0551_));
 NOR2_X1 _3421_ (.A1(prdata[6]),
    .A2(_1130_),
    .ZN(_1264_));
 AOI22_X1 _3422_ (.A1(\mem[14] [6]),
    .A2(net28),
    .B1(_1145_),
    .B2(\mem[1] [6]),
    .ZN(_1265_));
 NAND2_X1 _3423_ (.A1(\mem[9] [6]),
    .A2(net6),
    .ZN(_1266_));
 AOI22_X1 _3424_ (.A1(\mem[26] [6]),
    .A2(_1096_),
    .B1(net39),
    .B2(\mem[11] [6]),
    .ZN(_1267_));
 AOI22_X1 _3425_ (.A1(\mem[19] [6]),
    .A2(_1111_),
    .B1(_1140_),
    .B2(\mem[23] [6]),
    .ZN(_1268_));
 AOI22_X1 _3426_ (.A1(\mem[30] [6]),
    .A2(_1125_),
    .B1(_1143_),
    .B2(\mem[29] [6]),
    .ZN(_1269_));
 AOI22_X1 _3427_ (.A1(\mem[28] [6]),
    .A2(_1109_),
    .B1(_1146_),
    .B2(\mem[25] [6]),
    .ZN(_1270_));
 AND4_X1 _3428_ (.A1(_1267_),
    .A2(_1268_),
    .A3(_1269_),
    .A4(_1270_),
    .ZN(_1271_));
 AOI222_X2 _3429_ (.A1(\mem[15] [6]),
    .A2(net13),
    .B1(_1113_),
    .B2(\mem[24] [6]),
    .C1(net33),
    .C2(\mem[13] [6]),
    .ZN(_1272_));
 NAND2_X1 _3430_ (.A1(_1266_),
    .A2(_1272_),
    .ZN(_1273_));
 AOI222_X1 _3431_ (.A1(\mem[2] [6]),
    .A2(_1120_),
    .B1(_1123_),
    .B2(\mem[21] [6]),
    .C1(net44),
    .C2(\mem[3] [6]),
    .ZN(_1274_));
 AOI22_X1 _3432_ (.A1(\mem[5] [6]),
    .A2(_1138_),
    .B1(_1147_),
    .B2(\mem[6] [6]),
    .ZN(_1275_));
 NAND3_X1 _3433_ (.A1(_1265_),
    .A2(_1274_),
    .A3(_1275_),
    .ZN(_1276_));
 AOI222_X1 _3434_ (.A1(\mem[17] [6]),
    .A2(net70),
    .B1(_1133_),
    .B2(\mem[0] [6]),
    .C1(net18),
    .C2(\mem[7] [6]),
    .ZN(_1277_));
 AOI221_X1 _3435_ (.A(net3),
    .B1(_1137_),
    .B2(\mem[4] [6]),
    .C1(net64),
    .C2(\mem[18] [6]),
    .ZN(_1278_));
 NAND2_X1 _3436_ (.A1(_1277_),
    .A2(_1278_),
    .ZN(_1279_));
 AOI22_X1 _3437_ (.A1(\mem[16] [6]),
    .A2(net10),
    .B1(_1128_),
    .B2(\mem[22] [6]),
    .ZN(_1280_));
 AOI22_X1 _3438_ (.A1(\mem[20] [6]),
    .A2(_1118_),
    .B1(net22),
    .B2(\mem[8] [6]),
    .ZN(_1281_));
 AOI22_X1 _3439_ (.A1(\mem[12] [6]),
    .A2(_1077_),
    .B1(_1135_),
    .B2(\mem[10] [6]),
    .ZN(_1282_));
 AOI22_X1 _3440_ (.A1(\mem[31] [6]),
    .A2(_1101_),
    .B1(net66),
    .B2(\mem[27] [6]),
    .ZN(_1283_));
 NAND4_X1 _3441_ (.A1(_1280_),
    .A2(_1281_),
    .A3(_1282_),
    .A4(_1283_),
    .ZN(_1284_));
 NOR4_X1 _3442_ (.A1(_1273_),
    .A2(_1276_),
    .A3(_1279_),
    .A4(_1284_),
    .ZN(_1285_));
 AOI21_X1 _3443_ (.A(_1264_),
    .B1(_1271_),
    .B2(_1285_),
    .ZN(_0552_));
 NOR2_X1 _3444_ (.A1(prdata[7]),
    .A2(_1130_),
    .ZN(_1286_));
 AOI22_X1 _3445_ (.A1(\mem[18] [7]),
    .A2(net64),
    .B1(net36),
    .B2(\mem[23] [7]),
    .ZN(_1287_));
 AOI22_X1 _3446_ (.A1(\mem[0] [7]),
    .A2(net45),
    .B1(net44),
    .B2(\mem[3] [7]),
    .ZN(_1288_));
 AOI22_X1 _3447_ (.A1(\mem[5] [7]),
    .A2(_1138_),
    .B1(net24),
    .B2(\mem[1] [7]),
    .ZN(_1289_));
 AOI22_X1 _3448_ (.A1(\mem[25] [7]),
    .A2(_1146_),
    .B1(_1147_),
    .B2(\mem[6] [7]),
    .ZN(_1290_));
 AND4_X1 _3449_ (.A1(_1287_),
    .A2(_1288_),
    .A3(_1289_),
    .A4(_1290_),
    .ZN(_1291_));
 AOI222_X2 _3450_ (.A1(\mem[13] [7]),
    .A2(net32),
    .B1(net27),
    .B2(\mem[14] [7]),
    .C1(net21),
    .C2(\mem[8] [7]),
    .ZN(_1292_));
 AOI222_X1 _3451_ (.A1(\mem[20] [7]),
    .A2(net55),
    .B1(_1128_),
    .B2(\mem[22] [7]),
    .C1(net17),
    .C2(\mem[7] [7]),
    .ZN(_1293_));
 AOI22_X1 _3452_ (.A1(\mem[26] [7]),
    .A2(_1096_),
    .B1(net66),
    .B2(\mem[27] [7]),
    .ZN(_1294_));
 AOI222_X1 _3453_ (.A1(\mem[16] [7]),
    .A2(net11),
    .B1(net6),
    .B2(\mem[9] [7]),
    .C1(_1135_),
    .C2(\mem[10] [7]),
    .ZN(_1295_));
 NAND4_X1 _3454_ (.A1(_1292_),
    .A2(_1293_),
    .A3(_1294_),
    .A4(_1295_),
    .ZN(_1296_));
 AOI222_X1 _3455_ (.A1(\mem[12] [7]),
    .A2(_1077_),
    .B1(net12),
    .B2(\mem[15] [7]),
    .C1(_1139_),
    .C2(\mem[11] [7]),
    .ZN(_1297_));
 AOI221_X1 _3456_ (.A(net4),
    .B1(net47),
    .B2(\mem[30] [7]),
    .C1(\mem[31] [7]),
    .C2(_1101_),
    .ZN(_1298_));
 NAND2_X1 _3457_ (.A1(_1297_),
    .A2(_1298_),
    .ZN(_1299_));
 AOI22_X1 _3458_ (.A1(\mem[28] [7]),
    .A2(net61),
    .B1(net40),
    .B2(\mem[4] [7]),
    .ZN(_1300_));
 AOI22_X1 _3459_ (.A1(\mem[19] [7]),
    .A2(net60),
    .B1(net51),
    .B2(\mem[2] [7]),
    .ZN(_1301_));
 AOI22_X1 _3460_ (.A1(\mem[17] [7]),
    .A2(net68),
    .B1(_1123_),
    .B2(\mem[21] [7]),
    .ZN(_1302_));
 AOI22_X1 _3461_ (.A1(\mem[24] [7]),
    .A2(net57),
    .B1(_1143_),
    .B2(\mem[29] [7]),
    .ZN(_1303_));
 NAND4_X1 _3462_ (.A1(_1300_),
    .A2(_1301_),
    .A3(_1302_),
    .A4(_1303_),
    .ZN(_1304_));
 NOR3_X1 _3463_ (.A1(_1296_),
    .A2(_1299_),
    .A3(_1304_),
    .ZN(_1305_));
 AOI21_X1 _3464_ (.A(_1286_),
    .B1(_1291_),
    .B2(_1305_),
    .ZN(_0553_));
 NOR2_X1 _3465_ (.A1(prdata[8]),
    .A2(_1130_),
    .ZN(_1306_));
 NAND2_X1 _3466_ (.A1(\mem[19] [8]),
    .A2(_1111_),
    .ZN(_1307_));
 AOI222_X1 _3467_ (.A1(\mem[16] [8]),
    .A2(_1099_),
    .B1(_1128_),
    .B2(\mem[22] [8]),
    .C1(_1140_),
    .C2(\mem[23] [8]),
    .ZN(_1308_));
 AOI22_X1 _3468_ (.A1(\mem[17] [8]),
    .A2(_1103_),
    .B1(_1107_),
    .B2(\mem[18] [8]),
    .ZN(_1309_));
 AOI222_X1 _3469_ (.A1(\mem[12] [8]),
    .A2(_1077_),
    .B1(net13),
    .B2(\mem[15] [8]),
    .C1(net39),
    .C2(\mem[11] [8]),
    .ZN(_1310_));
 AND2_X1 _3470_ (.A1(_1309_),
    .A2(_1310_),
    .ZN(_1311_));
 AOI222_X1 _3471_ (.A1(\mem[5] [8]),
    .A2(_1138_),
    .B1(_1147_),
    .B2(\mem[6] [8]),
    .C1(_1145_),
    .C2(\mem[1] [8]),
    .ZN(_1312_));
 AOI22_X1 _3472_ (.A1(\mem[20] [8]),
    .A2(net55),
    .B1(net18),
    .B2(\mem[7] [8]),
    .ZN(_1313_));
 NAND2_X1 _3473_ (.A1(_1312_),
    .A2(_1313_),
    .ZN(_1314_));
 AOI221_X1 _3474_ (.A(net4),
    .B1(_1133_),
    .B2(\mem[0] [8]),
    .C1(net44),
    .C2(\mem[3] [8]),
    .ZN(_1315_));
 AOI222_X1 _3475_ (.A1(\mem[26] [8]),
    .A2(_1096_),
    .B1(_1120_),
    .B2(\mem[2] [8]),
    .C1(_1137_),
    .C2(\mem[4] [8]),
    .ZN(_1316_));
 NAND2_X1 _3476_ (.A1(_1315_),
    .A2(_1316_),
    .ZN(_1317_));
 AOI222_X1 _3477_ (.A1(\mem[31] [8]),
    .A2(net8),
    .B1(_1125_),
    .B2(\mem[30] [8]),
    .C1(_1143_),
    .C2(\mem[29] [8]),
    .ZN(_1318_));
 AOI22_X1 _3478_ (.A1(\mem[28] [8]),
    .A2(_1109_),
    .B1(_1146_),
    .B2(\mem[25] [8]),
    .ZN(_1319_));
 AOI22_X1 _3479_ (.A1(\mem[27] [8]),
    .A2(net66),
    .B1(_1113_),
    .B2(\mem[24] [8]),
    .ZN(_1320_));
 NAND3_X1 _3480_ (.A1(_1318_),
    .A2(_1319_),
    .A3(_1320_),
    .ZN(_1321_));
 AOI222_X2 _3481_ (.A1(\mem[13] [8]),
    .A2(_1141_),
    .B1(_1142_),
    .B2(\mem[14] [8]),
    .C1(_1148_),
    .C2(\mem[8] [8]),
    .ZN(_1322_));
 AOI222_X1 _3482_ (.A1(\mem[9] [8]),
    .A2(net6),
    .B1(_1123_),
    .B2(\mem[21] [8]),
    .C1(_1135_),
    .C2(\mem[10] [8]),
    .ZN(_1323_));
 NAND4_X1 _3483_ (.A1(_1307_),
    .A2(_1308_),
    .A3(_1322_),
    .A4(_1323_),
    .ZN(_1324_));
 NOR4_X1 _3484_ (.A1(_1314_),
    .A2(_1317_),
    .A3(_1321_),
    .A4(_1324_),
    .ZN(_1325_));
 AOI21_X1 _3485_ (.A(_1306_),
    .B1(_1311_),
    .B2(_1325_),
    .ZN(_0554_));
 NOR2_X1 _3486_ (.A1(prdata[9]),
    .A2(_1130_),
    .ZN(_1326_));
 AOI22_X1 _3487_ (.A1(\mem[18] [9]),
    .A2(_1107_),
    .B1(_1140_),
    .B2(\mem[23] [9]),
    .ZN(_1327_));
 AOI22_X1 _3488_ (.A1(\mem[11] [9]),
    .A2(net39),
    .B1(net33),
    .B2(\mem[13] [9]),
    .ZN(_1328_));
 AOI22_X1 _3489_ (.A1(\mem[12] [9]),
    .A2(net14),
    .B1(net6),
    .B2(\mem[9] [9]),
    .ZN(_1329_));
 AOI22_X1 _3490_ (.A1(\mem[14] [9]),
    .A2(net30),
    .B1(_1146_),
    .B2(\mem[25] [9]),
    .ZN(_1330_));
 AND4_X1 _3491_ (.A1(_1327_),
    .A2(_1328_),
    .A3(_1329_),
    .A4(_1330_),
    .ZN(_1331_));
 AOI222_X1 _3492_ (.A1(\mem[4] [9]),
    .A2(net42),
    .B1(_1147_),
    .B2(\mem[6] [9]),
    .C1(net24),
    .C2(\mem[1] [9]),
    .ZN(_1332_));
 AOI222_X2 _3493_ (.A1(\mem[20] [9]),
    .A2(_1118_),
    .B1(_1128_),
    .B2(\mem[22] [9]),
    .C1(net22),
    .C2(\mem[8] [9]),
    .ZN(_1333_));
 AOI22_X1 _3494_ (.A1(\mem[26] [9]),
    .A2(_1096_),
    .B1(_1105_),
    .B2(\mem[27] [9]),
    .ZN(_1334_));
 AOI222_X1 _3495_ (.A1(\mem[16] [9]),
    .A2(net10),
    .B1(net52),
    .B2(\mem[2] [9]),
    .C1(_1134_),
    .C2(\mem[3] [9]),
    .ZN(_1335_));
 NAND4_X1 _3496_ (.A1(_1332_),
    .A2(_1333_),
    .A3(_1334_),
    .A4(_1335_),
    .ZN(_1336_));
 AOI222_X1 _3497_ (.A1(\mem[0] [9]),
    .A2(net46),
    .B1(_1138_),
    .B2(\mem[5] [9]),
    .C1(\mem[7] [9]),
    .C2(_1149_),
    .ZN(_1337_));
 AOI221_X1 _3498_ (.A(net3),
    .B1(net49),
    .B2(\mem[30] [9]),
    .C1(\mem[31] [9]),
    .C2(net8),
    .ZN(_1338_));
 NAND2_X1 _3499_ (.A1(_1337_),
    .A2(_1338_),
    .ZN(_1339_));
 AOI22_X1 _3500_ (.A1(\mem[28] [9]),
    .A2(_1109_),
    .B1(_1135_),
    .B2(\mem[10] [9]),
    .ZN(_1340_));
 AOI22_X1 _3501_ (.A1(\mem[15] [9]),
    .A2(net13),
    .B1(_1111_),
    .B2(\mem[19] [9]),
    .ZN(_1341_));
 AOI22_X1 _3502_ (.A1(\mem[17] [9]),
    .A2(_1103_),
    .B1(_1123_),
    .B2(\mem[21] [9]),
    .ZN(_1342_));
 AOI22_X1 _3503_ (.A1(\mem[24] [9]),
    .A2(_1113_),
    .B1(net25),
    .B2(\mem[29] [9]),
    .ZN(_1343_));
 NAND4_X1 _3504_ (.A1(_1340_),
    .A2(_1341_),
    .A3(_1342_),
    .A4(_1343_),
    .ZN(_1344_));
 NOR3_X1 _3505_ (.A1(_1336_),
    .A2(_1339_),
    .A3(_1344_),
    .ZN(_1345_));
 AOI21_X1 _3506_ (.A(_1326_),
    .B1(_1331_),
    .B2(_1345_),
    .ZN(_0555_));
 NOR2_X1 _3507_ (.A1(prdata[10]),
    .A2(_1130_),
    .ZN(_1346_));
 AOI22_X1 _3508_ (.A1(\mem[16] [10]),
    .A2(net9),
    .B1(net50),
    .B2(\mem[2] [10]),
    .ZN(_1347_));
 AOI22_X1 _3509_ (.A1(\mem[18] [10]),
    .A2(net65),
    .B1(net59),
    .B2(\mem[19] [10]),
    .ZN(_1348_));
 AOI222_X1 _3510_ (.A1(\mem[15] [10]),
    .A2(net12),
    .B1(net53),
    .B2(\mem[20] [10]),
    .C1(net37),
    .C2(\mem[11] [10]),
    .ZN(_1349_));
 AOI221_X1 _3511_ (.A(_1131_),
    .B1(net35),
    .B2(\mem[23] [10]),
    .C1(net31),
    .C2(\mem[13] [10]),
    .ZN(_1350_));
 NAND2_X1 _3512_ (.A1(_1349_),
    .A2(_1350_),
    .ZN(_1351_));
 AOI22_X1 _3513_ (.A1(\mem[21] [10]),
    .A2(_1123_),
    .B1(_1128_),
    .B2(\mem[22] [10]),
    .ZN(_1352_));
 AOI22_X1 _3514_ (.A1(\mem[12] [10]),
    .A2(net15),
    .B1(net28),
    .B2(\mem[14] [10]),
    .ZN(_1353_));
 AOI22_X1 _3515_ (.A1(\mem[4] [10]),
    .A2(net41),
    .B1(_1146_),
    .B2(\mem[25] [10]),
    .ZN(_1354_));
 NAND4_X1 _3516_ (.A1(_1347_),
    .A2(_1352_),
    .A3(_1353_),
    .A4(_1354_),
    .ZN(_1355_));
 NOR2_X1 _3517_ (.A1(_1351_),
    .A2(_1355_),
    .ZN(_1356_));
 AOI222_X1 _3518_ (.A1(\mem[1] [10]),
    .A2(net23),
    .B1(net16),
    .B2(\mem[7] [10]),
    .C1(\mem[5] [10]),
    .C2(_1138_),
    .ZN(_1357_));
 AOI222_X1 _3519_ (.A1(\mem[28] [10]),
    .A2(net62),
    .B1(net56),
    .B2(\mem[24] [10]),
    .C1(_1147_),
    .C2(\mem[6] [10]),
    .ZN(_1358_));
 AOI222_X1 _3520_ (.A1(\mem[31] [10]),
    .A2(net7),
    .B1(net48),
    .B2(\mem[30] [10]),
    .C1(net26),
    .C2(\mem[29] [10]),
    .ZN(_1359_));
 NAND4_X1 _3521_ (.A1(_1348_),
    .A2(_1357_),
    .A3(_1358_),
    .A4(_1359_),
    .ZN(_1360_));
 AOI22_X1 _3522_ (.A1(\mem[0] [10]),
    .A2(net46),
    .B1(net43),
    .B2(\mem[3] [10]),
    .ZN(_1361_));
 AOI22_X1 _3523_ (.A1(\mem[17] [10]),
    .A2(net69),
    .B1(net19),
    .B2(\mem[8] [10]),
    .ZN(_1362_));
 AOI22_X1 _3524_ (.A1(\mem[9] [10]),
    .A2(net5),
    .B1(_1135_),
    .B2(\mem[10] [10]),
    .ZN(_1363_));
 AOI22_X1 _3525_ (.A1(\mem[26] [10]),
    .A2(_1096_),
    .B1(net67),
    .B2(\mem[27] [10]),
    .ZN(_1364_));
 NAND4_X1 _3526_ (.A1(_1361_),
    .A2(_1362_),
    .A3(_1363_),
    .A4(_1364_),
    .ZN(_1365_));
 NOR2_X1 _3527_ (.A1(_1360_),
    .A2(_1365_),
    .ZN(_1366_));
 AOI21_X1 _3528_ (.A(_1346_),
    .B1(_1356_),
    .B2(_1366_),
    .ZN(_0556_));
 NOR2_X1 _3529_ (.A1(prdata[11]),
    .A2(_1130_),
    .ZN(_1367_));
 AOI22_X1 _3530_ (.A1(\mem[18] [11]),
    .A2(net65),
    .B1(_1140_),
    .B2(\mem[23] [11]),
    .ZN(_1368_));
 AOI22_X1 _3531_ (.A1(\mem[27] [11]),
    .A2(net67),
    .B1(net58),
    .B2(\mem[24] [11]),
    .ZN(_1369_));
 AOI22_X1 _3532_ (.A1(\mem[29] [11]),
    .A2(net25),
    .B1(_1146_),
    .B2(\mem[25] [11]),
    .ZN(_1370_));
 AOI22_X1 _3533_ (.A1(\mem[12] [11]),
    .A2(net14),
    .B1(net8),
    .B2(\mem[31] [11]),
    .ZN(_1371_));
 AND4_X1 _3534_ (.A1(_1368_),
    .A2(_1369_),
    .A3(_1370_),
    .A4(_1371_),
    .ZN(_1372_));
 AOI222_X1 _3535_ (.A1(\mem[10] [11]),
    .A2(_1135_),
    .B1(_1147_),
    .B2(\mem[6] [11]),
    .C1(_1149_),
    .C2(\mem[7] [11]),
    .ZN(_1373_));
 AOI22_X1 _3536_ (.A1(\mem[15] [11]),
    .A2(_1093_),
    .B1(net20),
    .B2(\mem[8] [11]),
    .ZN(_1374_));
 AOI222_X1 _3537_ (.A1(\mem[20] [11]),
    .A2(net54),
    .B1(net48),
    .B2(\mem[30] [11]),
    .C1(_1128_),
    .C2(\mem[22] [11]),
    .ZN(_1375_));
 AOI222_X2 _3538_ (.A1(\mem[16] [11]),
    .A2(net10),
    .B1(_1138_),
    .B2(\mem[5] [11]),
    .C1(net30),
    .C2(\mem[14] [11]),
    .ZN(_1376_));
 NAND4_X1 _3539_ (.A1(_1373_),
    .A2(_1374_),
    .A3(_1375_),
    .A4(_1376_),
    .ZN(_1377_));
 AOI222_X1 _3540_ (.A1(\mem[0] [11]),
    .A2(net46),
    .B1(net42),
    .B2(\mem[4] [11]),
    .C1(net38),
    .C2(\mem[11] [11]),
    .ZN(_1378_));
 AOI221_X1 _3541_ (.A(net3),
    .B1(_1134_),
    .B2(\mem[3] [11]),
    .C1(net52),
    .C2(\mem[2] [11]),
    .ZN(_1379_));
 NAND2_X1 _3542_ (.A1(_1378_),
    .A2(_1379_),
    .ZN(_1380_));
 AOI22_X1 _3543_ (.A1(\mem[28] [11]),
    .A2(_1109_),
    .B1(net33),
    .B2(\mem[13] [11]),
    .ZN(_1381_));
 AOI22_X1 _3544_ (.A1(\mem[26] [11]),
    .A2(_1096_),
    .B1(_1111_),
    .B2(\mem[19] [11]),
    .ZN(_1382_));
 AOI22_X1 _3545_ (.A1(\mem[17] [11]),
    .A2(_1103_),
    .B1(_1123_),
    .B2(\mem[21] [11]),
    .ZN(_1383_));
 AOI22_X1 _3546_ (.A1(\mem[9] [11]),
    .A2(net6),
    .B1(_1145_),
    .B2(\mem[1] [11]),
    .ZN(_1384_));
 NAND4_X1 _3547_ (.A1(_1381_),
    .A2(_1382_),
    .A3(_1383_),
    .A4(_1384_),
    .ZN(_1385_));
 NOR3_X1 _3548_ (.A1(_1377_),
    .A2(_1380_),
    .A3(_1385_),
    .ZN(_1386_));
 AOI21_X1 _3549_ (.A(_1367_),
    .B1(_1372_),
    .B2(_1386_),
    .ZN(_0557_));
 AOI222_X1 _3550_ (.A1(\mem[5] [12]),
    .A2(_1138_),
    .B1(_1147_),
    .B2(\mem[6] [12]),
    .C1(_1145_),
    .C2(\mem[1] [12]),
    .ZN(_1387_));
 AOI22_X1 _3551_ (.A1(\mem[26] [12]),
    .A2(_1096_),
    .B1(net44),
    .B2(\mem[3] [12]),
    .ZN(_1388_));
 AOI222_X2 _3552_ (.A1(\mem[20] [12]),
    .A2(_1118_),
    .B1(_1128_),
    .B2(\mem[22] [12]),
    .C1(net27),
    .C2(\mem[14] [12]),
    .ZN(_1389_));
 AOI222_X1 _3553_ (.A1(\mem[16] [12]),
    .A2(net11),
    .B1(net66),
    .B2(\mem[27] [12]),
    .C1(_1120_),
    .C2(\mem[2] [12]),
    .ZN(_1390_));
 NAND4_X1 _3554_ (.A1(_1387_),
    .A2(_1388_),
    .A3(_1389_),
    .A4(_1390_),
    .ZN(_1391_));
 AOI22_X1 _3555_ (.A1(\mem[28] [12]),
    .A2(net61),
    .B1(net40),
    .B2(\mem[4] [12]),
    .ZN(_1392_));
 AOI222_X1 _3556_ (.A1(\mem[31] [12]),
    .A2(net7),
    .B1(net45),
    .B2(\mem[0] [12]),
    .C1(net18),
    .C2(\mem[7] [12]),
    .ZN(_1393_));
 AOI221_X1 _3557_ (.A(net3),
    .B1(net38),
    .B2(\mem[11] [12]),
    .C1(_1077_),
    .C2(\mem[12] [12]),
    .ZN(_1394_));
 AOI222_X1 _3558_ (.A1(\mem[15] [12]),
    .A2(_1093_),
    .B1(net57),
    .B2(\mem[24] [12]),
    .C1(_1135_),
    .C2(\mem[10] [12]),
    .ZN(_1395_));
 NAND4_X1 _3559_ (.A1(_1392_),
    .A2(_1393_),
    .A3(_1394_),
    .A4(_1395_),
    .ZN(_1396_));
 AOI22_X1 _3560_ (.A1(\mem[18] [12]),
    .A2(net64),
    .B1(net60),
    .B2(\mem[19] [12]),
    .ZN(_1397_));
 AOI222_X1 _3561_ (.A1(\mem[17] [12]),
    .A2(net68),
    .B1(_1123_),
    .B2(\mem[21] [12]),
    .C1(net36),
    .C2(\mem[23] [12]),
    .ZN(_1398_));
 AOI222_X2 _3562_ (.A1(\mem[9] [12]),
    .A2(_1116_),
    .B1(net32),
    .B2(\mem[13] [12]),
    .C1(net21),
    .C2(\mem[8] [12]),
    .ZN(_1399_));
 NAND3_X1 _3563_ (.A1(_1397_),
    .A2(_1398_),
    .A3(_1399_),
    .ZN(_1400_));
 AOI222_X1 _3564_ (.A1(\mem[30] [12]),
    .A2(_1125_),
    .B1(_1143_),
    .B2(\mem[29] [12]),
    .C1(_1146_),
    .C2(\mem[25] [12]),
    .ZN(_1401_));
 INV_X1 _3565_ (.A(_1401_),
    .ZN(_1402_));
 NOR4_X1 _3566_ (.A1(_1391_),
    .A2(_1396_),
    .A3(_1400_),
    .A4(_1402_),
    .ZN(_1403_));
 AOI21_X1 _3567_ (.A(_1403_),
    .B1(net4),
    .B2(_1062_),
    .ZN(_0558_));
 NOR2_X1 _3568_ (.A1(prdata[13]),
    .A2(_1130_),
    .ZN(_1404_));
 AOI22_X1 _3569_ (.A1(\mem[26] [13]),
    .A2(_1096_),
    .B1(net28),
    .B2(\mem[14] [13]),
    .ZN(_1405_));
 AOI22_X1 _3570_ (.A1(\mem[22] [13]),
    .A2(_1128_),
    .B1(net36),
    .B2(\mem[23] [13]),
    .ZN(_1406_));
 AOI22_X1 _3571_ (.A1(\mem[28] [13]),
    .A2(net61),
    .B1(_1146_),
    .B2(\mem[25] [13]),
    .ZN(_1407_));
 AOI22_X1 _3572_ (.A1(\mem[31] [13]),
    .A2(net7),
    .B1(net26),
    .B2(\mem[29] [13]),
    .ZN(_1408_));
 AND4_X1 _3573_ (.A1(_1405_),
    .A2(_1406_),
    .A3(_1407_),
    .A4(_1408_),
    .ZN(_1409_));
 AOI222_X1 _3574_ (.A1(\mem[9] [13]),
    .A2(net5),
    .B1(net51),
    .B2(\mem[2] [13]),
    .C1(net24),
    .C2(\mem[1] [13]),
    .ZN(_1410_));
 AOI22_X1 _3575_ (.A1(\mem[10] [13]),
    .A2(_1135_),
    .B1(net34),
    .B2(\mem[13] [13]),
    .ZN(_1411_));
 NAND2_X1 _3576_ (.A1(_1410_),
    .A2(_1411_),
    .ZN(_1412_));
 AOI222_X2 _3577_ (.A1(\mem[21] [13]),
    .A2(_1123_),
    .B1(_1138_),
    .B2(\mem[5] [13]),
    .C1(net21),
    .C2(\mem[8] [13]),
    .ZN(_1413_));
 AOI222_X1 _3578_ (.A1(\mem[4] [13]),
    .A2(net40),
    .B1(_1147_),
    .B2(\mem[6] [13]),
    .C1(net17),
    .C2(\mem[7] [13]),
    .ZN(_1414_));
 NAND2_X1 _3579_ (.A1(_1413_),
    .A2(_1414_),
    .ZN(_1415_));
 AOI222_X1 _3580_ (.A1(\mem[17] [13]),
    .A2(net68),
    .B1(net45),
    .B2(\mem[0] [13]),
    .C1(net37),
    .C2(\mem[11] [13]),
    .ZN(_1416_));
 AOI221_X1 _3581_ (.A(net4),
    .B1(net60),
    .B2(\mem[19] [13]),
    .C1(\mem[18] [13]),
    .C2(net63),
    .ZN(_1417_));
 NAND2_X1 _3582_ (.A1(_1416_),
    .A2(_1417_),
    .ZN(_1418_));
 AOI22_X1 _3583_ (.A1(\mem[16] [13]),
    .A2(net11),
    .B1(net53),
    .B2(\mem[20] [13]),
    .ZN(_1419_));
 AOI22_X1 _3584_ (.A1(\mem[12] [13]),
    .A2(net15),
    .B1(net12),
    .B2(\mem[15] [13]),
    .ZN(_1420_));
 AOI22_X1 _3585_ (.A1(\mem[27] [13]),
    .A2(_1105_),
    .B1(net56),
    .B2(\mem[24] [13]),
    .ZN(_1421_));
 AOI22_X1 _3586_ (.A1(\mem[30] [13]),
    .A2(net47),
    .B1(net44),
    .B2(\mem[3] [13]),
    .ZN(_1422_));
 NAND4_X1 _3587_ (.A1(_1419_),
    .A2(_1420_),
    .A3(_1421_),
    .A4(_1422_),
    .ZN(_1423_));
 NOR4_X1 _3588_ (.A1(_1412_),
    .A2(_1415_),
    .A3(_1418_),
    .A4(_1423_),
    .ZN(_1424_));
 AOI21_X1 _3589_ (.A(_1404_),
    .B1(_1409_),
    .B2(_1424_),
    .ZN(_0559_));
 NOR2_X1 _3590_ (.A1(prdata[14]),
    .A2(_1130_),
    .ZN(_1425_));
 AOI22_X1 _3591_ (.A1(\mem[18] [14]),
    .A2(net64),
    .B1(net60),
    .B2(\mem[19] [14]),
    .ZN(_1426_));
 AOI22_X1 _3592_ (.A1(\mem[20] [14]),
    .A2(net55),
    .B1(net45),
    .B2(\mem[0] [14]),
    .ZN(_1427_));
 AOI22_X1 _3593_ (.A1(\mem[5] [14]),
    .A2(_1138_),
    .B1(net24),
    .B2(\mem[1] [14]),
    .ZN(_1428_));
 AOI22_X1 _3594_ (.A1(\mem[12] [14]),
    .A2(net15),
    .B1(net40),
    .B2(\mem[4] [14]),
    .ZN(_1429_));
 AOI22_X1 _3595_ (.A1(\mem[11] [14]),
    .A2(net37),
    .B1(net36),
    .B2(\mem[23] [14]),
    .ZN(_1430_));
 AND4_X1 _3596_ (.A1(_1427_),
    .A2(_1428_),
    .A3(_1429_),
    .A4(_1430_),
    .ZN(_1431_));
 AOI222_X2 _3597_ (.A1(\mem[15] [14]),
    .A2(net12),
    .B1(net6),
    .B2(\mem[9] [14]),
    .C1(net32),
    .C2(\mem[13] [14]),
    .ZN(_1432_));
 AOI222_X2 _3598_ (.A1(\mem[28] [14]),
    .A2(net61),
    .B1(net56),
    .B2(\mem[24] [14]),
    .C1(net27),
    .C2(\mem[14] [14]),
    .ZN(_1433_));
 AOI222_X1 _3599_ (.A1(\mem[31] [14]),
    .A2(_1101_),
    .B1(net47),
    .B2(\mem[30] [14]),
    .C1(_1143_),
    .C2(\mem[29] [14]),
    .ZN(_1434_));
 NAND4_X1 _3600_ (.A1(_1426_),
    .A2(_1432_),
    .A3(_1433_),
    .A4(_1434_),
    .ZN(_1435_));
 AOI222_X1 _3601_ (.A1(\mem[17] [14]),
    .A2(net68),
    .B1(_1123_),
    .B2(\mem[21] [14]),
    .C1(_1128_),
    .C2(\mem[22] [14]),
    .ZN(_1436_));
 AOI221_X1 _3602_ (.A(net4),
    .B1(_1147_),
    .B2(\mem[6] [14]),
    .C1(net11),
    .C2(\mem[16] [14]),
    .ZN(_1437_));
 NAND2_X1 _3603_ (.A1(_1436_),
    .A2(_1437_),
    .ZN(_1438_));
 AOI22_X1 _3604_ (.A1(\mem[2] [14]),
    .A2(net51),
    .B1(net44),
    .B2(\mem[3] [14]),
    .ZN(_1439_));
 AOI22_X1 _3605_ (.A1(\mem[27] [14]),
    .A2(net66),
    .B1(net17),
    .B2(\mem[7] [14]),
    .ZN(_1440_));
 AOI22_X1 _3606_ (.A1(\mem[26] [14]),
    .A2(_1096_),
    .B1(_1146_),
    .B2(\mem[25] [14]),
    .ZN(_1441_));
 AOI22_X1 _3607_ (.A1(\mem[10] [14]),
    .A2(_1135_),
    .B1(net21),
    .B2(\mem[8] [14]),
    .ZN(_1442_));
 NAND4_X1 _3608_ (.A1(_1439_),
    .A2(_1440_),
    .A3(_1441_),
    .A4(_1442_),
    .ZN(_1443_));
 NOR3_X1 _3609_ (.A1(_1435_),
    .A2(_1438_),
    .A3(_1443_),
    .ZN(_1444_));
 AOI21_X1 _3610_ (.A(_1425_),
    .B1(_1431_),
    .B2(_1444_),
    .ZN(_0560_));
 NOR2_X1 _3611_ (.A1(prdata[15]),
    .A2(_1130_),
    .ZN(_1445_));
 AOI22_X1 _3612_ (.A1(\mem[1] [15]),
    .A2(net24),
    .B1(_1147_),
    .B2(\mem[6] [15]),
    .ZN(_1446_));
 NAND2_X1 _3613_ (.A1(\mem[15] [15]),
    .A2(net12),
    .ZN(_1447_));
 AOI22_X1 _3614_ (.A1(\mem[12] [15]),
    .A2(net15),
    .B1(_1096_),
    .B2(\mem[26] [15]),
    .ZN(_1448_));
 AOI22_X1 _3615_ (.A1(\mem[22] [15]),
    .A2(_1128_),
    .B1(net36),
    .B2(\mem[23] [15]),
    .ZN(_1449_));
 AOI22_X1 _3616_ (.A1(\mem[28] [15]),
    .A2(net61),
    .B1(_1146_),
    .B2(\mem[25] [15]),
    .ZN(_1450_));
 AOI22_X1 _3617_ (.A1(\mem[31] [15]),
    .A2(net7),
    .B1(net26),
    .B2(\mem[29] [15]),
    .ZN(_1451_));
 AND4_X1 _3618_ (.A1(_1448_),
    .A2(_1449_),
    .A3(_1450_),
    .A4(_1451_),
    .ZN(_1452_));
 AOI222_X2 _3619_ (.A1(\mem[9] [15]),
    .A2(net6),
    .B1(net32),
    .B2(\mem[13] [15]),
    .C1(net27),
    .C2(\mem[14] [15]),
    .ZN(_1453_));
 NAND2_X1 _3620_ (.A1(_1447_),
    .A2(_1453_),
    .ZN(_1454_));
 AOI222_X1 _3621_ (.A1(\mem[21] [15]),
    .A2(_1123_),
    .B1(net44),
    .B2(\mem[3] [15]),
    .C1(net41),
    .C2(\mem[4] [15]),
    .ZN(_1455_));
 AOI22_X1 _3622_ (.A1(\mem[2] [15]),
    .A2(net51),
    .B1(_1138_),
    .B2(\mem[5] [15]),
    .ZN(_1456_));
 NAND3_X1 _3623_ (.A1(_1446_),
    .A2(_1455_),
    .A3(_1456_),
    .ZN(_1457_));
 AOI222_X1 _3624_ (.A1(\mem[17] [15]),
    .A2(net68),
    .B1(net45),
    .B2(\mem[0] [15]),
    .C1(net17),
    .C2(\mem[7] [15]),
    .ZN(_1458_));
 AOI221_X1 _3625_ (.A(net4),
    .B1(net60),
    .B2(\mem[19] [15]),
    .C1(\mem[18] [15]),
    .C2(net64),
    .ZN(_1459_));
 NAND2_X1 _3626_ (.A1(_1458_),
    .A2(_1459_),
    .ZN(_1460_));
 AOI22_X1 _3627_ (.A1(\mem[16] [15]),
    .A2(net9),
    .B1(net55),
    .B2(\mem[20] [15]),
    .ZN(_1461_));
 AOI22_X1 _3628_ (.A1(\mem[11] [15]),
    .A2(net37),
    .B1(net21),
    .B2(\mem[8] [15]),
    .ZN(_1462_));
 AOI22_X1 _3629_ (.A1(\mem[27] [15]),
    .A2(net66),
    .B1(net56),
    .B2(\mem[24] [15]),
    .ZN(_1463_));
 AOI22_X1 _3630_ (.A1(\mem[30] [15]),
    .A2(net47),
    .B1(_1135_),
    .B2(\mem[10] [15]),
    .ZN(_1464_));
 NAND4_X1 _3631_ (.A1(_1461_),
    .A2(_1462_),
    .A3(_1463_),
    .A4(_1464_),
    .ZN(_1465_));
 NOR4_X1 _3632_ (.A1(_1454_),
    .A2(_1457_),
    .A3(_1460_),
    .A4(_1465_),
    .ZN(_1466_));
 AOI21_X1 _3633_ (.A(_1445_),
    .B1(_1452_),
    .B2(_1466_),
    .ZN(_0561_));
 NOR2_X1 _3634_ (.A1(prdata[16]),
    .A2(_1130_),
    .ZN(_1467_));
 AOI22_X1 _3635_ (.A1(\mem[16] [16]),
    .A2(net9),
    .B1(net54),
    .B2(\mem[20] [16]),
    .ZN(_1468_));
 AOI222_X1 _3636_ (.A1(\mem[1] [16]),
    .A2(net23),
    .B1(net18),
    .B2(\mem[7] [16]),
    .C1(\mem[4] [16]),
    .C2(net42),
    .ZN(_1469_));
 AOI221_X1 _3637_ (.A(net3),
    .B1(_1147_),
    .B2(\mem[6] [16]),
    .C1(net60),
    .C2(\mem[19] [16]),
    .ZN(_1470_));
 AOI22_X1 _3638_ (.A1(\mem[0] [16]),
    .A2(net46),
    .B1(net43),
    .B2(\mem[3] [16]),
    .ZN(_1471_));
 AOI22_X1 _3639_ (.A1(\mem[27] [16]),
    .A2(_1105_),
    .B1(net57),
    .B2(\mem[24] [16]),
    .ZN(_1472_));
 AOI22_X1 _3640_ (.A1(\mem[2] [16]),
    .A2(net52),
    .B1(net48),
    .B2(\mem[30] [16]),
    .ZN(_1473_));
 AND4_X1 _3641_ (.A1(_1468_),
    .A2(_1471_),
    .A3(_1472_),
    .A4(_1473_),
    .ZN(_1474_));
 AND3_X1 _3642_ (.A1(_1469_),
    .A2(_1470_),
    .A3(_1474_),
    .ZN(_1475_));
 AOI222_X2 _3643_ (.A1(\mem[12] [16]),
    .A2(_1077_),
    .B1(net29),
    .B2(\mem[14] [16]),
    .C1(net20),
    .C2(\mem[8] [16]),
    .ZN(_1476_));
 INV_X1 _3644_ (.A(_1476_),
    .ZN(_1477_));
 AOI22_X1 _3645_ (.A1(\mem[9] [16]),
    .A2(net5),
    .B1(_1123_),
    .B2(\mem[21] [16]),
    .ZN(_1478_));
 AOI22_X1 _3646_ (.A1(\mem[10] [16]),
    .A2(_1135_),
    .B1(net34),
    .B2(\mem[13] [16]),
    .ZN(_1479_));
 AOI22_X1 _3647_ (.A1(\mem[17] [16]),
    .A2(net69),
    .B1(net65),
    .B2(\mem[18] [16]),
    .ZN(_1480_));
 AOI22_X1 _3648_ (.A1(\mem[15] [16]),
    .A2(_1093_),
    .B1(net38),
    .B2(\mem[11] [16]),
    .ZN(_1481_));
 NAND4_X1 _3649_ (.A1(_1478_),
    .A2(_1479_),
    .A3(_1480_),
    .A4(_1481_),
    .ZN(_1482_));
 AOI22_X1 _3650_ (.A1(\mem[22] [16]),
    .A2(_1128_),
    .B1(net35),
    .B2(\mem[23] [16]),
    .ZN(_1483_));
 AOI22_X1 _3651_ (.A1(\mem[26] [16]),
    .A2(_1096_),
    .B1(_1138_),
    .B2(\mem[5] [16]),
    .ZN(_1484_));
 AOI22_X1 _3652_ (.A1(\mem[31] [16]),
    .A2(net8),
    .B1(net62),
    .B2(\mem[28] [16]),
    .ZN(_1485_));
 AOI22_X1 _3653_ (.A1(\mem[29] [16]),
    .A2(net25),
    .B1(_1146_),
    .B2(\mem[25] [16]),
    .ZN(_1486_));
 NAND4_X1 _3654_ (.A1(_1483_),
    .A2(_1484_),
    .A3(_1485_),
    .A4(_1486_),
    .ZN(_1487_));
 NOR3_X1 _3655_ (.A1(_1477_),
    .A2(_1482_),
    .A3(_1487_),
    .ZN(_1488_));
 AOI21_X1 _3656_ (.A(_1467_),
    .B1(_1475_),
    .B2(_1488_),
    .ZN(_0562_));
 NOR2_X1 _3657_ (.A1(prdata[17]),
    .A2(_1130_),
    .ZN(_1489_));
 AOI22_X1 _3658_ (.A1(\mem[2] [17]),
    .A2(net52),
    .B1(net43),
    .B2(\mem[3] [17]),
    .ZN(_1490_));
 AOI222_X2 _3659_ (.A1(\mem[16] [17]),
    .A2(net9),
    .B1(net70),
    .B2(\mem[17] [17]),
    .C1(_1123_),
    .C2(\mem[21] [17]),
    .ZN(_1491_));
 AOI221_X1 _3660_ (.A(net3),
    .B1(_1147_),
    .B2(\mem[6] [17]),
    .C1(net54),
    .C2(\mem[20] [17]),
    .ZN(_1492_));
 NAND2_X1 _3661_ (.A1(_1491_),
    .A2(_1492_),
    .ZN(_1493_));
 AOI22_X1 _3662_ (.A1(\mem[27] [17]),
    .A2(_1105_),
    .B1(net16),
    .B2(\mem[7] [17]),
    .ZN(_1494_));
 AOI22_X1 _3663_ (.A1(\mem[26] [17]),
    .A2(_1096_),
    .B1(_1146_),
    .B2(\mem[25] [17]),
    .ZN(_1495_));
 AOI22_X1 _3664_ (.A1(\mem[10] [17]),
    .A2(_1135_),
    .B1(net19),
    .B2(\mem[8] [17]),
    .ZN(_1496_));
 NAND4_X1 _3665_ (.A1(_1490_),
    .A2(_1494_),
    .A3(_1495_),
    .A4(_1496_),
    .ZN(_1497_));
 NOR2_X1 _3666_ (.A1(_1493_),
    .A2(_1497_),
    .ZN(_1498_));
 AOI22_X1 _3667_ (.A1(\mem[18] [17]),
    .A2(net63),
    .B1(net59),
    .B2(\mem[19] [17]),
    .ZN(_1499_));
 AOI222_X2 _3668_ (.A1(\mem[9] [17]),
    .A2(net5),
    .B1(net31),
    .B2(\mem[13] [17]),
    .C1(net29),
    .C2(\mem[14] [17]),
    .ZN(_1500_));
 AOI222_X1 _3669_ (.A1(\mem[15] [17]),
    .A2(_1093_),
    .B1(net62),
    .B2(\mem[28] [17]),
    .C1(net57),
    .C2(\mem[24] [17]),
    .ZN(_1501_));
 AOI222_X1 _3670_ (.A1(\mem[31] [17]),
    .A2(net8),
    .B1(net48),
    .B2(\mem[30] [17]),
    .C1(net25),
    .C2(\mem[29] [17]),
    .ZN(_1502_));
 NAND4_X1 _3671_ (.A1(_1499_),
    .A2(_1500_),
    .A3(_1501_),
    .A4(_1502_),
    .ZN(_1503_));
 AOI22_X1 _3672_ (.A1(\mem[4] [17]),
    .A2(net42),
    .B1(net23),
    .B2(\mem[1] [17]),
    .ZN(_1504_));
 AOI22_X1 _3673_ (.A1(\mem[22] [17]),
    .A2(_1128_),
    .B1(net46),
    .B2(\mem[0] [17]),
    .ZN(_1505_));
 AOI22_X1 _3674_ (.A1(\mem[12] [17]),
    .A2(_1077_),
    .B1(net35),
    .B2(\mem[23] [17]),
    .ZN(_1506_));
 AOI22_X1 _3675_ (.A1(\mem[5] [17]),
    .A2(_1138_),
    .B1(net38),
    .B2(\mem[11] [17]),
    .ZN(_1507_));
 NAND4_X1 _3676_ (.A1(_1504_),
    .A2(_1505_),
    .A3(_1506_),
    .A4(_1507_),
    .ZN(_1508_));
 NOR2_X1 _3677_ (.A1(_1503_),
    .A2(_1508_),
    .ZN(_1509_));
 AOI21_X1 _3678_ (.A(_1489_),
    .B1(_1498_),
    .B2(_1509_),
    .ZN(_0563_));
 NOR2_X1 _3679_ (.A1(prdata[18]),
    .A2(_1130_),
    .ZN(_1510_));
 AOI22_X1 _3680_ (.A1(\mem[2] [18]),
    .A2(net52),
    .B1(_1123_),
    .B2(\mem[21] [18]),
    .ZN(_1511_));
 AOI222_X1 _3681_ (.A1(\mem[26] [18]),
    .A2(_1096_),
    .B1(_1111_),
    .B2(\mem[19] [18]),
    .C1(net35),
    .C2(\mem[23] [18]),
    .ZN(_1512_));
 AOI221_X1 _3682_ (.A(_1131_),
    .B1(net65),
    .B2(\mem[18] [18]),
    .C1(\mem[27] [18]),
    .C2(net67),
    .ZN(_1513_));
 NAND2_X1 _3683_ (.A1(_1512_),
    .A2(_1513_),
    .ZN(_1514_));
 AOI22_X1 _3684_ (.A1(\mem[0] [18]),
    .A2(net46),
    .B1(_1145_),
    .B2(\mem[1] [18]),
    .ZN(_1515_));
 AOI22_X1 _3685_ (.A1(\mem[20] [18]),
    .A2(net54),
    .B1(net25),
    .B2(\mem[29] [18]),
    .ZN(_1516_));
 AOI22_X1 _3686_ (.A1(\mem[9] [18]),
    .A2(net5),
    .B1(_1134_),
    .B2(\mem[3] [18]),
    .ZN(_1517_));
 NAND4_X1 _3687_ (.A1(_1511_),
    .A2(_1515_),
    .A3(_1516_),
    .A4(_1517_),
    .ZN(_1518_));
 NOR2_X1 _3688_ (.A1(_1514_),
    .A2(_1518_),
    .ZN(_1519_));
 AOI222_X1 _3689_ (.A1(\mem[15] [18]),
    .A2(net13),
    .B1(_1135_),
    .B2(\mem[10] [18]),
    .C1(net39),
    .C2(\mem[11] [18]),
    .ZN(_1520_));
 AOI22_X1 _3690_ (.A1(\mem[28] [18]),
    .A2(_1109_),
    .B1(net22),
    .B2(\mem[8] [18]),
    .ZN(_1521_));
 AOI222_X2 _3691_ (.A1(\mem[12] [18]),
    .A2(net14),
    .B1(_1138_),
    .B2(\mem[5] [18]),
    .C1(net30),
    .C2(\mem[14] [18]),
    .ZN(_1522_));
 AOI222_X1 _3692_ (.A1(\mem[31] [18]),
    .A2(net8),
    .B1(net58),
    .B2(\mem[24] [18]),
    .C1(net49),
    .C2(\mem[30] [18]),
    .ZN(_1523_));
 NAND4_X1 _3693_ (.A1(_1520_),
    .A2(_1521_),
    .A3(_1522_),
    .A4(_1523_),
    .ZN(_1524_));
 AOI22_X1 _3694_ (.A1(\mem[22] [18]),
    .A2(_1128_),
    .B1(_1146_),
    .B2(\mem[25] [18]),
    .ZN(_1525_));
 AOI22_X1 _3695_ (.A1(\mem[16] [18]),
    .A2(net10),
    .B1(_1147_),
    .B2(\mem[6] [18]),
    .ZN(_1526_));
 AOI22_X1 _3696_ (.A1(\mem[17] [18]),
    .A2(net69),
    .B1(_1149_),
    .B2(\mem[7] [18]),
    .ZN(_1527_));
 AOI22_X1 _3697_ (.A1(\mem[4] [18]),
    .A2(net42),
    .B1(net33),
    .B2(\mem[13] [18]),
    .ZN(_1528_));
 NAND4_X1 _3698_ (.A1(_1525_),
    .A2(_1526_),
    .A3(_1527_),
    .A4(_1528_),
    .ZN(_1529_));
 NOR2_X1 _3699_ (.A1(_1524_),
    .A2(_1529_),
    .ZN(_1530_));
 AOI21_X1 _3700_ (.A(_1510_),
    .B1(_1519_),
    .B2(_1530_),
    .ZN(_0564_));
 AOI222_X2 _3701_ (.A1(\mem[13] [19]),
    .A2(net33),
    .B1(net30),
    .B2(\mem[14] [19]),
    .C1(net22),
    .C2(\mem[8] [19]),
    .ZN(_1531_));
 AOI222_X1 _3702_ (.A1(\mem[20] [19]),
    .A2(net54),
    .B1(_1128_),
    .B2(\mem[22] [19]),
    .C1(_1147_),
    .C2(\mem[6] [19]),
    .ZN(_1532_));
 AOI22_X1 _3703_ (.A1(\mem[26] [19]),
    .A2(_1096_),
    .B1(net67),
    .B2(\mem[27] [19]),
    .ZN(_1533_));
 AOI222_X1 _3704_ (.A1(\mem[16] [19]),
    .A2(_1099_),
    .B1(net6),
    .B2(\mem[9] [19]),
    .C1(_1135_),
    .C2(\mem[10] [19]),
    .ZN(_1534_));
 NAND4_X1 _3705_ (.A1(_1531_),
    .A2(_1532_),
    .A3(_1533_),
    .A4(_1534_),
    .ZN(_1535_));
 AOI22_X1 _3706_ (.A1(\mem[12] [19]),
    .A2(net14),
    .B1(net8),
    .B2(\mem[31] [19]),
    .ZN(_1536_));
 AOI222_X1 _3707_ (.A1(\mem[15] [19]),
    .A2(net13),
    .B1(_1109_),
    .B2(\mem[28] [19]),
    .C1(net39),
    .C2(\mem[11] [19]),
    .ZN(_1537_));
 AOI221_X1 _3708_ (.A(net3),
    .B1(net46),
    .B2(\mem[0] [19]),
    .C1(_1134_),
    .C2(\mem[3] [19]),
    .ZN(_1538_));
 AOI222_X1 _3709_ (.A1(\mem[24] [19]),
    .A2(net58),
    .B1(net52),
    .B2(\mem[2] [19]),
    .C1(_1138_),
    .C2(\mem[5] [19]),
    .ZN(_1539_));
 NAND4_X1 _3710_ (.A1(_1536_),
    .A2(_1537_),
    .A3(_1538_),
    .A4(_1539_),
    .ZN(_1540_));
 AOI22_X1 _3711_ (.A1(\mem[18] [19]),
    .A2(_1107_),
    .B1(_1111_),
    .B2(\mem[19] [19]),
    .ZN(_1541_));
 AOI222_X1 _3712_ (.A1(\mem[17] [19]),
    .A2(_1103_),
    .B1(_1123_),
    .B2(\mem[21] [19]),
    .C1(_1140_),
    .C2(\mem[23] [19]),
    .ZN(_1542_));
 AOI222_X1 _3713_ (.A1(\mem[1] [19]),
    .A2(_1145_),
    .B1(_1149_),
    .B2(\mem[7] [19]),
    .C1(\mem[4] [19]),
    .C2(net42),
    .ZN(_1543_));
 NAND3_X1 _3714_ (.A1(_1541_),
    .A2(_1542_),
    .A3(_1543_),
    .ZN(_1544_));
 AOI222_X1 _3715_ (.A1(\mem[30] [19]),
    .A2(net49),
    .B1(net25),
    .B2(\mem[29] [19]),
    .C1(_1146_),
    .C2(\mem[25] [19]),
    .ZN(_1545_));
 INV_X1 _3716_ (.A(_1545_),
    .ZN(_1546_));
 NOR4_X1 _3717_ (.A1(_1535_),
    .A2(_1540_),
    .A3(_1544_),
    .A4(_1546_),
    .ZN(_1547_));
 AOI21_X1 _3718_ (.A(_1547_),
    .B1(net3),
    .B2(_1063_),
    .ZN(_0565_));
 AOI222_X1 _3719_ (.A1(\mem[10] [20]),
    .A2(_1135_),
    .B1(_1147_),
    .B2(\mem[6] [20]),
    .C1(net18),
    .C2(\mem[7] [20]),
    .ZN(_1548_));
 AOI22_X1 _3720_ (.A1(\mem[9] [20]),
    .A2(net6),
    .B1(net27),
    .B2(\mem[14] [20]),
    .ZN(_1549_));
 AOI222_X1 _3721_ (.A1(\mem[20] [20]),
    .A2(net55),
    .B1(net47),
    .B2(\mem[30] [20]),
    .C1(_1128_),
    .C2(\mem[22] [20]),
    .ZN(_1550_));
 AOI222_X1 _3722_ (.A1(\mem[15] [20]),
    .A2(net13),
    .B1(_1099_),
    .B2(\mem[16] [20]),
    .C1(_1137_),
    .C2(\mem[4] [20]),
    .ZN(_1551_));
 NAND4_X1 _3723_ (.A1(_1548_),
    .A2(_1549_),
    .A3(_1550_),
    .A4(_1551_),
    .ZN(_1552_));
 AOI22_X1 _3724_ (.A1(\mem[0] [20]),
    .A2(_1133_),
    .B1(net44),
    .B2(\mem[3] [20]),
    .ZN(_1553_));
 AOI222_X1 _3725_ (.A1(\mem[2] [20]),
    .A2(_1120_),
    .B1(_1138_),
    .B2(\mem[5] [20]),
    .C1(_1139_),
    .C2(\mem[11] [20]),
    .ZN(_1554_));
 AOI221_X1 _3726_ (.A(net4),
    .B1(_1109_),
    .B2(\mem[28] [20]),
    .C1(\mem[27] [20]),
    .C2(net66),
    .ZN(_1555_));
 AOI222_X2 _3727_ (.A1(\mem[26] [20]),
    .A2(_1096_),
    .B1(_1101_),
    .B2(\mem[31] [20]),
    .C1(_1141_),
    .C2(\mem[13] [20]),
    .ZN(_1556_));
 NAND4_X1 _3728_ (.A1(_1553_),
    .A2(_1554_),
    .A3(_1555_),
    .A4(_1556_),
    .ZN(_1557_));
 AOI22_X1 _3729_ (.A1(\mem[18] [20]),
    .A2(net64),
    .B1(_1111_),
    .B2(\mem[19] [20]),
    .ZN(_1558_));
 AOI222_X1 _3730_ (.A1(\mem[17] [20]),
    .A2(_1103_),
    .B1(_1123_),
    .B2(\mem[21] [20]),
    .C1(_1140_),
    .C2(\mem[23] [20]),
    .ZN(_1559_));
 AOI222_X1 _3731_ (.A1(\mem[24] [20]),
    .A2(net57),
    .B1(_1143_),
    .B2(\mem[29] [20]),
    .C1(_1146_),
    .C2(\mem[25] [20]),
    .ZN(_1560_));
 NAND3_X1 _3732_ (.A1(_1558_),
    .A2(_1559_),
    .A3(_1560_),
    .ZN(_1561_));
 AOI222_X2 _3733_ (.A1(\mem[12] [20]),
    .A2(_1077_),
    .B1(_1145_),
    .B2(\mem[1] [20]),
    .C1(_1148_),
    .C2(\mem[8] [20]),
    .ZN(_1562_));
 INV_X1 _3734_ (.A(_1562_),
    .ZN(_1563_));
 NOR4_X1 _3735_ (.A1(_1552_),
    .A2(_1557_),
    .A3(_1561_),
    .A4(_1563_),
    .ZN(_1564_));
 AOI21_X1 _3736_ (.A(_1564_),
    .B1(net4),
    .B2(_1064_),
    .ZN(_0566_));
 NOR2_X1 _3737_ (.A1(prdata[21]),
    .A2(_1130_),
    .ZN(_1565_));
 AOI22_X1 _3738_ (.A1(\mem[4] [21]),
    .A2(net41),
    .B1(_1147_),
    .B2(\mem[6] [21]),
    .ZN(_1566_));
 AOI222_X1 _3739_ (.A1(\mem[20] [21]),
    .A2(net53),
    .B1(_1128_),
    .B2(\mem[22] [21]),
    .C1(_1135_),
    .C2(\mem[10] [21]),
    .ZN(_1567_));
 AOI221_X1 _3740_ (.A(_1131_),
    .B1(net48),
    .B2(\mem[30] [21]),
    .C1(\mem[28] [21]),
    .C2(net62),
    .ZN(_1568_));
 NAND2_X1 _3741_ (.A1(_1567_),
    .A2(_1568_),
    .ZN(_1569_));
 AOI22_X1 _3742_ (.A1(\mem[31] [21]),
    .A2(net7),
    .B1(net31),
    .B2(\mem[13] [21]),
    .ZN(_1570_));
 AOI22_X1 _3743_ (.A1(\mem[29] [21]),
    .A2(net26),
    .B1(net19),
    .B2(\mem[8] [21]),
    .ZN(_1571_));
 AOI22_X1 _3744_ (.A1(\mem[26] [21]),
    .A2(_1096_),
    .B1(net35),
    .B2(\mem[23] [21]),
    .ZN(_1572_));
 NAND4_X1 _3745_ (.A1(_1566_),
    .A2(_1570_),
    .A3(_1571_),
    .A4(_1572_),
    .ZN(_1573_));
 NOR2_X1 _3746_ (.A1(_1569_),
    .A2(_1573_),
    .ZN(_1574_));
 AOI222_X1 _3747_ (.A1(\mem[17] [21]),
    .A2(net69),
    .B1(_1123_),
    .B2(\mem[21] [21]),
    .C1(net43),
    .C2(\mem[3] [21]),
    .ZN(_1575_));
 AOI22_X1 _3748_ (.A1(\mem[19] [21]),
    .A2(net59),
    .B1(_1138_),
    .B2(\mem[5] [21]),
    .ZN(_1576_));
 AOI222_X2 _3749_ (.A1(\mem[12] [21]),
    .A2(net14),
    .B1(net5),
    .B2(\mem[9] [21]),
    .C1(net29),
    .C2(\mem[14] [21]),
    .ZN(_1577_));
 AOI222_X2 _3750_ (.A1(\mem[16] [21]),
    .A2(net10),
    .B1(net65),
    .B2(\mem[18] [21]),
    .C1(net46),
    .C2(\mem[0] [21]),
    .ZN(_1578_));
 NAND4_X1 _3751_ (.A1(_1575_),
    .A2(_1576_),
    .A3(_1577_),
    .A4(_1578_),
    .ZN(_1579_));
 AOI22_X1 _3752_ (.A1(\mem[27] [21]),
    .A2(net67),
    .B1(net16),
    .B2(\mem[7] [21]),
    .ZN(_1580_));
 AOI22_X1 _3753_ (.A1(\mem[15] [21]),
    .A2(_1093_),
    .B1(net38),
    .B2(\mem[11] [21]),
    .ZN(_1581_));
 AOI22_X1 _3754_ (.A1(\mem[2] [21]),
    .A2(net50),
    .B1(net23),
    .B2(\mem[1] [21]),
    .ZN(_1582_));
 AOI22_X1 _3755_ (.A1(\mem[24] [21]),
    .A2(net58),
    .B1(_1146_),
    .B2(\mem[25] [21]),
    .ZN(_1583_));
 NAND4_X1 _3756_ (.A1(_1580_),
    .A2(_1581_),
    .A3(_1582_),
    .A4(_1583_),
    .ZN(_1584_));
 NOR2_X1 _3757_ (.A1(_1579_),
    .A2(_1584_),
    .ZN(_1585_));
 AOI21_X1 _3758_ (.A(_1565_),
    .B1(_1574_),
    .B2(_1585_),
    .ZN(_0567_));
 NOR2_X1 _3759_ (.A1(prdata[22]),
    .A2(_1130_),
    .ZN(_1586_));
 AOI22_X1 _3760_ (.A1(\mem[20] [22]),
    .A2(net54),
    .B1(net50),
    .B2(\mem[2] [22]),
    .ZN(_1587_));
 AOI222_X2 _3761_ (.A1(\mem[15] [22]),
    .A2(net13),
    .B1(net39),
    .B2(\mem[11] [22]),
    .C1(net33),
    .C2(\mem[13] [22]),
    .ZN(_1588_));
 AOI221_X1 _3762_ (.A(net3),
    .B1(net35),
    .B2(\mem[23] [22]),
    .C1(_1128_),
    .C2(\mem[22] [22]),
    .ZN(_1589_));
 NAND2_X1 _3763_ (.A1(_1588_),
    .A2(_1589_),
    .ZN(_1590_));
 AOI22_X1 _3764_ (.A1(\mem[17] [22]),
    .A2(_1103_),
    .B1(_1123_),
    .B2(\mem[21] [22]),
    .ZN(_1591_));
 AOI22_X1 _3765_ (.A1(\mem[14] [22]),
    .A2(net30),
    .B1(net22),
    .B2(\mem[8] [22]),
    .ZN(_1592_));
 AOI22_X1 _3766_ (.A1(\mem[5] [22]),
    .A2(_1138_),
    .B1(_1146_),
    .B2(\mem[25] [22]),
    .ZN(_1593_));
 NAND4_X1 _3767_ (.A1(_1587_),
    .A2(_1591_),
    .A3(_1592_),
    .A4(_1593_),
    .ZN(_1594_));
 NOR2_X1 _3768_ (.A1(_1590_),
    .A2(_1594_),
    .ZN(_1595_));
 AOI222_X1 _3769_ (.A1(\mem[18] [22]),
    .A2(_1107_),
    .B1(_1109_),
    .B2(\mem[28] [22]),
    .C1(_1111_),
    .C2(\mem[19] [22]),
    .ZN(_1596_));
 AOI22_X1 _3770_ (.A1(\mem[24] [22]),
    .A2(net58),
    .B1(net25),
    .B2(\mem[29] [22]),
    .ZN(_1597_));
 AOI222_X1 _3771_ (.A1(\mem[1] [22]),
    .A2(_1145_),
    .B1(_1149_),
    .B2(\mem[7] [22]),
    .C1(\mem[4] [22]),
    .C2(net42),
    .ZN(_1598_));
 AOI222_X1 _3772_ (.A1(\mem[31] [22]),
    .A2(net8),
    .B1(net49),
    .B2(\mem[30] [22]),
    .C1(_1147_),
    .C2(\mem[6] [22]),
    .ZN(_1599_));
 NAND4_X1 _3773_ (.A1(_1596_),
    .A2(_1597_),
    .A3(_1598_),
    .A4(_1599_),
    .ZN(_1600_));
 AOI22_X1 _3774_ (.A1(\mem[0] [22]),
    .A2(net46),
    .B1(_1134_),
    .B2(\mem[3] [22]),
    .ZN(_1601_));
 AOI22_X1 _3775_ (.A1(\mem[12] [22]),
    .A2(net14),
    .B1(net10),
    .B2(\mem[16] [22]),
    .ZN(_1602_));
 AOI22_X1 _3776_ (.A1(\mem[9] [22]),
    .A2(net6),
    .B1(_1135_),
    .B2(\mem[10] [22]),
    .ZN(_1603_));
 AOI22_X1 _3777_ (.A1(\mem[26] [22]),
    .A2(_1096_),
    .B1(net67),
    .B2(\mem[27] [22]),
    .ZN(_1604_));
 NAND4_X1 _3778_ (.A1(_1601_),
    .A2(_1602_),
    .A3(_1603_),
    .A4(_1604_),
    .ZN(_1605_));
 NOR2_X1 _3779_ (.A1(_1600_),
    .A2(_1605_),
    .ZN(_1606_));
 AOI21_X1 _3780_ (.A(_1586_),
    .B1(_1595_),
    .B2(_1606_),
    .ZN(_0568_));
 NOR2_X1 _3781_ (.A1(prdata[23]),
    .A2(_1130_),
    .ZN(_1607_));
 AOI22_X1 _3782_ (.A1(\mem[18] [23]),
    .A2(net63),
    .B1(net36),
    .B2(\mem[23] [23]),
    .ZN(_1608_));
 AOI22_X1 _3783_ (.A1(\mem[27] [23]),
    .A2(_1105_),
    .B1(net61),
    .B2(\mem[28] [23]),
    .ZN(_1609_));
 AOI22_X1 _3784_ (.A1(\mem[24] [23]),
    .A2(net56),
    .B1(net26),
    .B2(\mem[29] [23]),
    .ZN(_1610_));
 AOI22_X1 _3785_ (.A1(\mem[12] [23]),
    .A2(net15),
    .B1(_1146_),
    .B2(\mem[25] [23]),
    .ZN(_1611_));
 AND4_X1 _3786_ (.A1(_1608_),
    .A2(_1609_),
    .A3(_1610_),
    .A4(_1611_),
    .ZN(_1612_));
 AOI222_X1 _3787_ (.A1(\mem[10] [23]),
    .A2(_1135_),
    .B1(_1147_),
    .B2(\mem[6] [23]),
    .C1(net17),
    .C2(\mem[7] [23]),
    .ZN(_1613_));
 AOI22_X1 _3788_ (.A1(\mem[9] [23]),
    .A2(_1116_),
    .B1(net28),
    .B2(\mem[14] [23]),
    .ZN(_1614_));
 AOI222_X1 _3789_ (.A1(\mem[20] [23]),
    .A2(net53),
    .B1(net47),
    .B2(\mem[30] [23]),
    .C1(_1128_),
    .C2(\mem[22] [23]),
    .ZN(_1615_));
 AOI222_X1 _3790_ (.A1(\mem[15] [23]),
    .A2(net12),
    .B1(net11),
    .B2(\mem[16] [23]),
    .C1(net40),
    .C2(\mem[4] [23]),
    .ZN(_1616_));
 NAND4_X1 _3791_ (.A1(_1613_),
    .A2(_1614_),
    .A3(_1615_),
    .A4(_1616_),
    .ZN(_1617_));
 AOI222_X1 _3792_ (.A1(\mem[0] [23]),
    .A2(net45),
    .B1(net37),
    .B2(\mem[11] [23]),
    .C1(_1138_),
    .C2(\mem[5] [23]),
    .ZN(_1618_));
 AOI221_X1 _3793_ (.A(net4),
    .B1(net44),
    .B2(\mem[3] [23]),
    .C1(net51),
    .C2(\mem[2] [23]),
    .ZN(_1619_));
 NAND2_X1 _3794_ (.A1(_1618_),
    .A2(_1619_),
    .ZN(_1620_));
 AOI22_X1 _3795_ (.A1(\mem[26] [23]),
    .A2(_1096_),
    .B1(net20),
    .B2(\mem[8] [23]),
    .ZN(_1621_));
 AOI22_X1 _3796_ (.A1(\mem[31] [23]),
    .A2(net7),
    .B1(net59),
    .B2(\mem[19] [23]),
    .ZN(_1622_));
 AOI22_X1 _3797_ (.A1(\mem[17] [23]),
    .A2(net68),
    .B1(_1123_),
    .B2(\mem[21] [23]),
    .ZN(_1623_));
 AOI22_X1 _3798_ (.A1(\mem[13] [23]),
    .A2(net34),
    .B1(net24),
    .B2(\mem[1] [23]),
    .ZN(_1624_));
 NAND4_X1 _3799_ (.A1(_1621_),
    .A2(_1622_),
    .A3(_1623_),
    .A4(_1624_),
    .ZN(_1625_));
 NOR3_X1 _3800_ (.A1(_1617_),
    .A2(_1620_),
    .A3(_1625_),
    .ZN(_1626_));
 AOI21_X1 _3801_ (.A(_1607_),
    .B1(_1612_),
    .B2(_1626_),
    .ZN(_0569_));
 NOR2_X1 _3802_ (.A1(prdata[24]),
    .A2(_1130_),
    .ZN(_1627_));
 AOI22_X1 _3803_ (.A1(\mem[2] [24]),
    .A2(net50),
    .B1(net43),
    .B2(\mem[3] [24]),
    .ZN(_1628_));
 AOI222_X1 _3804_ (.A1(\mem[17] [24]),
    .A2(net69),
    .B1(_1123_),
    .B2(\mem[21] [24]),
    .C1(_1128_),
    .C2(\mem[22] [24]),
    .ZN(_1629_));
 AOI221_X1 _3805_ (.A(_1131_),
    .B1(_1147_),
    .B2(\mem[6] [24]),
    .C1(net9),
    .C2(\mem[16] [24]),
    .ZN(_1630_));
 NAND2_X1 _3806_ (.A1(_1629_),
    .A2(_1630_),
    .ZN(_1631_));
 AOI22_X1 _3807_ (.A1(\mem[27] [24]),
    .A2(net67),
    .B1(net16),
    .B2(\mem[7] [24]),
    .ZN(_1632_));
 AOI22_X1 _3808_ (.A1(\mem[26] [24]),
    .A2(_1096_),
    .B1(_1146_),
    .B2(\mem[25] [24]),
    .ZN(_1633_));
 AOI22_X1 _3809_ (.A1(\mem[10] [24]),
    .A2(_1135_),
    .B1(net19),
    .B2(\mem[8] [24]),
    .ZN(_1634_));
 NAND4_X1 _3810_ (.A1(_1628_),
    .A2(_1632_),
    .A3(_1633_),
    .A4(_1634_),
    .ZN(_1635_));
 NOR2_X1 _3811_ (.A1(_1631_),
    .A2(_1635_),
    .ZN(_1636_));
 AOI22_X1 _3812_ (.A1(\mem[18] [24]),
    .A2(net65),
    .B1(net59),
    .B2(\mem[19] [24]),
    .ZN(_1637_));
 AOI222_X2 _3813_ (.A1(\mem[12] [24]),
    .A2(net14),
    .B1(net5),
    .B2(\mem[9] [24]),
    .C1(net29),
    .C2(\mem[14] [24]),
    .ZN(_1638_));
 AOI222_X2 _3814_ (.A1(\mem[15] [24]),
    .A2(_1093_),
    .B1(net62),
    .B2(\mem[28] [24]),
    .C1(net58),
    .C2(\mem[24] [24]),
    .ZN(_1639_));
 AOI222_X1 _3815_ (.A1(\mem[31] [24]),
    .A2(net7),
    .B1(net48),
    .B2(\mem[30] [24]),
    .C1(net26),
    .C2(\mem[29] [24]),
    .ZN(_1640_));
 NAND4_X1 _3816_ (.A1(_1637_),
    .A2(_1638_),
    .A3(_1639_),
    .A4(_1640_),
    .ZN(_1641_));
 AOI22_X1 _3817_ (.A1(\mem[5] [24]),
    .A2(_1138_),
    .B1(net23),
    .B2(\mem[1] [24]),
    .ZN(_1642_));
 AOI22_X1 _3818_ (.A1(\mem[20] [24]),
    .A2(net53),
    .B1(net46),
    .B2(\mem[0] [24]),
    .ZN(_1643_));
 AOI22_X1 _3819_ (.A1(\mem[4] [24]),
    .A2(net41),
    .B1(net31),
    .B2(\mem[13] [24]),
    .ZN(_1644_));
 AOI22_X1 _3820_ (.A1(\mem[11] [24]),
    .A2(net38),
    .B1(net35),
    .B2(\mem[23] [24]),
    .ZN(_1645_));
 NAND4_X1 _3821_ (.A1(_1642_),
    .A2(_1643_),
    .A3(_1644_),
    .A4(_1645_),
    .ZN(_1646_));
 NOR2_X1 _3822_ (.A1(_1641_),
    .A2(_1646_),
    .ZN(_1647_));
 AOI21_X1 _3823_ (.A(_1627_),
    .B1(_1636_),
    .B2(_1647_),
    .ZN(_0570_));
 AOI222_X2 _3824_ (.A1(\mem[13] [25]),
    .A2(net31),
    .B1(net29),
    .B2(\mem[14] [25]),
    .C1(net20),
    .C2(\mem[8] [25]),
    .ZN(_1648_));
 AOI222_X1 _3825_ (.A1(\mem[20] [25]),
    .A2(net53),
    .B1(_1128_),
    .B2(\mem[22] [25]),
    .C1(_1147_),
    .C2(\mem[6] [25]),
    .ZN(_1649_));
 AOI22_X1 _3826_ (.A1(\mem[26] [25]),
    .A2(_1096_),
    .B1(_1105_),
    .B2(\mem[27] [25]),
    .ZN(_1650_));
 AOI222_X1 _3827_ (.A1(\mem[16] [25]),
    .A2(net9),
    .B1(net5),
    .B2(\mem[9] [25]),
    .C1(_1135_),
    .C2(\mem[10] [25]),
    .ZN(_1651_));
 NAND4_X1 _3828_ (.A1(_1648_),
    .A2(_1649_),
    .A3(_1650_),
    .A4(_1651_),
    .ZN(_1652_));
 AOI22_X1 _3829_ (.A1(\mem[12] [25]),
    .A2(net15),
    .B1(net7),
    .B2(\mem[31] [25]),
    .ZN(_1653_));
 AOI222_X1 _3830_ (.A1(\mem[15] [25]),
    .A2(_1093_),
    .B1(net48),
    .B2(\mem[30] [25]),
    .C1(net37),
    .C2(\mem[11] [25]),
    .ZN(_1654_));
 AOI221_X1 _3831_ (.A(net3),
    .B1(net46),
    .B2(\mem[0] [25]),
    .C1(net43),
    .C2(\mem[3] [25]),
    .ZN(_1655_));
 AOI222_X1 _3832_ (.A1(\mem[28] [25]),
    .A2(net62),
    .B1(net52),
    .B2(\mem[2] [25]),
    .C1(net41),
    .C2(\mem[4] [25]),
    .ZN(_1656_));
 NAND4_X1 _3833_ (.A1(_1653_),
    .A2(_1654_),
    .A3(_1655_),
    .A4(_1656_),
    .ZN(_1657_));
 AOI22_X1 _3834_ (.A1(\mem[18] [25]),
    .A2(net63),
    .B1(net59),
    .B2(\mem[19] [25]),
    .ZN(_1658_));
 AOI222_X1 _3835_ (.A1(\mem[17] [25]),
    .A2(net70),
    .B1(_1123_),
    .B2(\mem[21] [25]),
    .C1(net36),
    .C2(\mem[23] [25]),
    .ZN(_1659_));
 AOI222_X1 _3836_ (.A1(\mem[1] [25]),
    .A2(net23),
    .B1(net18),
    .B2(\mem[7] [25]),
    .C1(\mem[5] [25]),
    .C2(_1138_),
    .ZN(_1660_));
 NAND3_X1 _3837_ (.A1(_1658_),
    .A2(_1659_),
    .A3(_1660_),
    .ZN(_1661_));
 AOI222_X1 _3838_ (.A1(\mem[24] [25]),
    .A2(net56),
    .B1(net26),
    .B2(\mem[29] [25]),
    .C1(_1146_),
    .C2(\mem[25] [25]),
    .ZN(_1662_));
 INV_X1 _3839_ (.A(_1662_),
    .ZN(_1663_));
 NOR4_X2 _3840_ (.A1(_1652_),
    .A2(_1657_),
    .A3(_1661_),
    .A4(_1663_),
    .ZN(_1664_));
 AOI21_X1 _3841_ (.A(_1664_),
    .B1(net3),
    .B2(_1065_),
    .ZN(_0571_));
 AOI222_X1 _3842_ (.A1(\mem[4] [26]),
    .A2(net42),
    .B1(_1147_),
    .B2(\mem[6] [26]),
    .C1(_1145_),
    .C2(\mem[1] [26]),
    .ZN(_1665_));
 AOI222_X2 _3843_ (.A1(\mem[20] [26]),
    .A2(net54),
    .B1(_1128_),
    .B2(\mem[22] [26]),
    .C1(net30),
    .C2(\mem[14] [26]),
    .ZN(_1666_));
 AOI22_X1 _3844_ (.A1(\mem[26] [26]),
    .A2(_1096_),
    .B1(net67),
    .B2(\mem[27] [26]),
    .ZN(_1667_));
 AOI222_X1 _3845_ (.A1(\mem[16] [26]),
    .A2(net10),
    .B1(net50),
    .B2(\mem[2] [26]),
    .C1(_1134_),
    .C2(\mem[3] [26]),
    .ZN(_1668_));
 NAND4_X1 _3846_ (.A1(_1665_),
    .A2(_1666_),
    .A3(_1667_),
    .A4(_1668_),
    .ZN(_1669_));
 AOI22_X1 _3847_ (.A1(\mem[31] [26]),
    .A2(net8),
    .B1(_1138_),
    .B2(\mem[5] [26]),
    .ZN(_1670_));
 AOI222_X1 _3848_ (.A1(\mem[30] [26]),
    .A2(net49),
    .B1(net46),
    .B2(\mem[0] [26]),
    .C1(_1149_),
    .C2(\mem[7] [26]),
    .ZN(_1671_));
 AOI221_X1 _3849_ (.A(_1131_),
    .B1(net39),
    .B2(\mem[11] [26]),
    .C1(net14),
    .C2(\mem[12] [26]),
    .ZN(_1672_));
 AOI222_X1 _3850_ (.A1(\mem[15] [26]),
    .A2(net13),
    .B1(_1109_),
    .B2(\mem[28] [26]),
    .C1(_1135_),
    .C2(\mem[10] [26]),
    .ZN(_1673_));
 NAND4_X1 _3851_ (.A1(_1670_),
    .A2(_1671_),
    .A3(_1672_),
    .A4(_1673_),
    .ZN(_1674_));
 AOI22_X1 _3852_ (.A1(\mem[18] [26]),
    .A2(_1107_),
    .B1(_1111_),
    .B2(\mem[19] [26]),
    .ZN(_1675_));
 AOI222_X1 _3853_ (.A1(\mem[17] [26]),
    .A2(_1103_),
    .B1(_1123_),
    .B2(\mem[21] [26]),
    .C1(net35),
    .C2(\mem[23] [26]),
    .ZN(_1676_));
 AOI222_X2 _3854_ (.A1(\mem[9] [26]),
    .A2(net6),
    .B1(net33),
    .B2(\mem[13] [26]),
    .C1(net22),
    .C2(\mem[8] [26]),
    .ZN(_1677_));
 NAND3_X1 _3855_ (.A1(_1675_),
    .A2(_1676_),
    .A3(_1677_),
    .ZN(_1678_));
 AOI222_X1 _3856_ (.A1(\mem[24] [26]),
    .A2(net58),
    .B1(net25),
    .B2(\mem[29] [26]),
    .C1(_1146_),
    .C2(\mem[25] [26]),
    .ZN(_1679_));
 INV_X1 _3857_ (.A(_1679_),
    .ZN(_1680_));
 NOR4_X1 _3858_ (.A1(_1669_),
    .A2(_1674_),
    .A3(_1678_),
    .A4(_1680_),
    .ZN(_1681_));
 AOI21_X1 _3859_ (.A(_1681_),
    .B1(_1131_),
    .B2(_1066_),
    .ZN(_0572_));
 AOI222_X2 _3860_ (.A1(\mem[12] [27]),
    .A2(_1077_),
    .B1(_1142_),
    .B2(\mem[14] [27]),
    .C1(_1148_),
    .C2(\mem[8] [27]),
    .ZN(_1682_));
 AOI222_X1 _3861_ (.A1(\mem[20] [27]),
    .A2(net55),
    .B1(_1128_),
    .B2(\mem[22] [27]),
    .C1(_1147_),
    .C2(\mem[6] [27]),
    .ZN(_1683_));
 AOI22_X1 _3862_ (.A1(\mem[26] [27]),
    .A2(_1096_),
    .B1(net66),
    .B2(\mem[27] [27]),
    .ZN(_1684_));
 AOI222_X1 _3863_ (.A1(\mem[16] [27]),
    .A2(_1099_),
    .B1(net6),
    .B2(\mem[9] [27]),
    .C1(_1135_),
    .C2(\mem[10] [27]),
    .ZN(_1685_));
 NAND4_X1 _3864_ (.A1(_1682_),
    .A2(_1683_),
    .A3(_1684_),
    .A4(_1685_),
    .ZN(_1686_));
 AOI22_X1 _3865_ (.A1(\mem[28] [27]),
    .A2(_1109_),
    .B1(_1141_),
    .B2(\mem[13] [27]),
    .ZN(_1687_));
 AOI222_X1 _3866_ (.A1(\mem[15] [27]),
    .A2(net13),
    .B1(net8),
    .B2(\mem[31] [27]),
    .C1(net39),
    .C2(\mem[11] [27]),
    .ZN(_1688_));
 AOI221_X1 _3867_ (.A(net3),
    .B1(_1133_),
    .B2(\mem[0] [27]),
    .C1(net44),
    .C2(\mem[3] [27]),
    .ZN(_1689_));
 AOI222_X2 _3868_ (.A1(\mem[24] [27]),
    .A2(net57),
    .B1(_1120_),
    .B2(\mem[2] [27]),
    .C1(_1137_),
    .C2(\mem[4] [27]),
    .ZN(_1690_));
 NAND4_X1 _3869_ (.A1(_1687_),
    .A2(_1688_),
    .A3(_1689_),
    .A4(_1690_),
    .ZN(_1691_));
 AOI22_X1 _3870_ (.A1(\mem[18] [27]),
    .A2(_1107_),
    .B1(_1111_),
    .B2(\mem[19] [27]),
    .ZN(_1692_));
 AOI222_X1 _3871_ (.A1(\mem[17] [27]),
    .A2(_1103_),
    .B1(_1123_),
    .B2(\mem[21] [27]),
    .C1(_1140_),
    .C2(\mem[23] [27]),
    .ZN(_1693_));
 AOI222_X1 _3872_ (.A1(\mem[1] [27]),
    .A2(_1145_),
    .B1(net18),
    .B2(\mem[7] [27]),
    .C1(\mem[5] [27]),
    .C2(_1138_),
    .ZN(_1694_));
 NAND3_X1 _3873_ (.A1(_1692_),
    .A2(_1693_),
    .A3(_1694_),
    .ZN(_1695_));
 AOI222_X1 _3874_ (.A1(\mem[30] [27]),
    .A2(_1125_),
    .B1(_1143_),
    .B2(\mem[29] [27]),
    .C1(_1146_),
    .C2(\mem[25] [27]),
    .ZN(_1696_));
 INV_X1 _3875_ (.A(_1696_),
    .ZN(_1697_));
 NOR4_X1 _3876_ (.A1(_1686_),
    .A2(_1691_),
    .A3(_1695_),
    .A4(_1697_),
    .ZN(_1698_));
 AOI21_X1 _3877_ (.A(_1698_),
    .B1(net3),
    .B2(_1067_),
    .ZN(_0573_));
 NOR2_X1 _3878_ (.A1(prdata[28]),
    .A2(_1130_),
    .ZN(_1699_));
 AOI22_X1 _3879_ (.A1(\mem[18] [28]),
    .A2(net63),
    .B1(net36),
    .B2(\mem[23] [28]),
    .ZN(_1700_));
 AOI22_X1 _3880_ (.A1(\mem[11] [28]),
    .A2(net37),
    .B1(net21),
    .B2(\mem[8] [28]),
    .ZN(_1701_));
 AOI22_X1 _3881_ (.A1(\mem[9] [28]),
    .A2(net5),
    .B1(net34),
    .B2(\mem[13] [28]),
    .ZN(_1702_));
 AOI22_X1 _3882_ (.A1(\mem[15] [28]),
    .A2(net12),
    .B1(_1146_),
    .B2(\mem[25] [28]),
    .ZN(_1703_));
 AND4_X1 _3883_ (.A1(_1700_),
    .A2(_1701_),
    .A3(_1702_),
    .A4(_1703_),
    .ZN(_1704_));
 AOI222_X1 _3884_ (.A1(\mem[4] [28]),
    .A2(net41),
    .B1(_1147_),
    .B2(\mem[6] [28]),
    .C1(net24),
    .C2(\mem[1] [28]),
    .ZN(_1705_));
 AOI222_X2 _3885_ (.A1(\mem[20] [28]),
    .A2(net55),
    .B1(_1128_),
    .B2(\mem[22] [28]),
    .C1(net28),
    .C2(\mem[14] [28]),
    .ZN(_1706_));
 AOI22_X1 _3886_ (.A1(\mem[26] [28]),
    .A2(_1096_),
    .B1(net66),
    .B2(\mem[27] [28]),
    .ZN(_1707_));
 AOI222_X1 _3887_ (.A1(\mem[16] [28]),
    .A2(net9),
    .B1(net51),
    .B2(\mem[2] [28]),
    .C1(net44),
    .C2(\mem[3] [28]),
    .ZN(_1708_));
 NAND4_X1 _3888_ (.A1(_1705_),
    .A2(_1706_),
    .A3(_1707_),
    .A4(_1708_),
    .ZN(_1709_));
 AOI222_X1 _3889_ (.A1(\mem[0] [28]),
    .A2(net45),
    .B1(_1138_),
    .B2(\mem[5] [28]),
    .C1(\mem[7] [28]),
    .C2(net17),
    .ZN(_1710_));
 AOI221_X1 _3890_ (.A(net4),
    .B1(net47),
    .B2(\mem[30] [28]),
    .C1(\mem[31] [28]),
    .C2(net7),
    .ZN(_1711_));
 NAND2_X1 _3891_ (.A1(_1710_),
    .A2(_1711_),
    .ZN(_1712_));
 AOI22_X1 _3892_ (.A1(\mem[12] [28]),
    .A2(net15),
    .B1(net61),
    .B2(\mem[28] [28]),
    .ZN(_1713_));
 AOI22_X1 _3893_ (.A1(\mem[19] [28]),
    .A2(net60),
    .B1(_1135_),
    .B2(\mem[10] [28]),
    .ZN(_1714_));
 AOI22_X1 _3894_ (.A1(\mem[17] [28]),
    .A2(net68),
    .B1(_1123_),
    .B2(\mem[21] [28]),
    .ZN(_1715_));
 AOI22_X1 _3895_ (.A1(\mem[24] [28]),
    .A2(net56),
    .B1(net26),
    .B2(\mem[29] [28]),
    .ZN(_1716_));
 NAND4_X1 _3896_ (.A1(_1713_),
    .A2(_1714_),
    .A3(_1715_),
    .A4(_1716_),
    .ZN(_1717_));
 NOR3_X1 _3897_ (.A1(_1709_),
    .A2(_1712_),
    .A3(_1717_),
    .ZN(_1718_));
 AOI21_X1 _3898_ (.A(_1699_),
    .B1(_1704_),
    .B2(_1718_),
    .ZN(_0574_));
 NOR2_X1 _3899_ (.A1(prdata[29]),
    .A2(_1130_),
    .ZN(_1719_));
 AOI222_X1 _3900_ (.A1(\mem[20] [29]),
    .A2(_1118_),
    .B1(_1128_),
    .B2(\mem[22] [29]),
    .C1(_1135_),
    .C2(\mem[10] [29]),
    .ZN(_1720_));
 INV_X1 _3901_ (.A(_1720_),
    .ZN(_1721_));
 AOI222_X2 _3902_ (.A1(\mem[9] [29]),
    .A2(net6),
    .B1(net32),
    .B2(\mem[13] [29]),
    .C1(net27),
    .C2(\mem[14] [29]),
    .ZN(_1722_));
 AOI221_X1 _3903_ (.A(net4),
    .B1(net57),
    .B2(\mem[24] [29]),
    .C1(\mem[27] [29]),
    .C2(net66),
    .ZN(_1723_));
 AOI22_X1 _3904_ (.A1(\mem[5] [29]),
    .A2(_1138_),
    .B1(net17),
    .B2(\mem[7] [29]),
    .ZN(_1724_));
 AOI22_X1 _3905_ (.A1(\mem[26] [29]),
    .A2(_1096_),
    .B1(_1147_),
    .B2(\mem[6] [29]),
    .ZN(_1725_));
 NAND3_X1 _3906_ (.A1(_1723_),
    .A2(_1724_),
    .A3(_1725_),
    .ZN(_1726_));
 AOI211_X2 _3907_ (.A(_1721_),
    .B(_1726_),
    .C1(\mem[30] [29]),
    .C2(net47),
    .ZN(_1727_));
 AOI22_X1 _3908_ (.A1(\mem[12] [29]),
    .A2(_1077_),
    .B1(net13),
    .B2(\mem[15] [29]),
    .ZN(_1728_));
 INV_X1 _3909_ (.A(_1728_),
    .ZN(_1729_));
 AOI22_X1 _3910_ (.A1(\mem[11] [29]),
    .A2(_1139_),
    .B1(net21),
    .B2(\mem[8] [29]),
    .ZN(_1730_));
 AOI222_X1 _3911_ (.A1(\mem[31] [29]),
    .A2(_1101_),
    .B1(_1143_),
    .B2(\mem[29] [29]),
    .C1(_1146_),
    .C2(\mem[25] [29]),
    .ZN(_1731_));
 AOI222_X1 _3912_ (.A1(\mem[28] [29]),
    .A2(net61),
    .B1(net51),
    .B2(\mem[2] [29]),
    .C1(_1145_),
    .C2(\mem[1] [29]),
    .ZN(_1732_));
 NAND3_X1 _3913_ (.A1(_1730_),
    .A2(_1731_),
    .A3(_1732_),
    .ZN(_1733_));
 AOI222_X1 _3914_ (.A1(\mem[17] [29]),
    .A2(_1103_),
    .B1(_1123_),
    .B2(\mem[21] [29]),
    .C1(_1140_),
    .C2(\mem[23] [29]),
    .ZN(_1734_));
 AOI222_X1 _3915_ (.A1(\mem[16] [29]),
    .A2(net11),
    .B1(net44),
    .B2(\mem[3] [29]),
    .C1(_1137_),
    .C2(\mem[4] [29]),
    .ZN(_1735_));
 AOI222_X1 _3916_ (.A1(\mem[18] [29]),
    .A2(net64),
    .B1(net60),
    .B2(\mem[19] [29]),
    .C1(_1133_),
    .C2(\mem[0] [29]),
    .ZN(_1736_));
 NAND4_X1 _3917_ (.A1(_1722_),
    .A2(_1734_),
    .A3(_1735_),
    .A4(_1736_),
    .ZN(_1737_));
 NOR3_X1 _3918_ (.A1(_1729_),
    .A2(_1733_),
    .A3(_1737_),
    .ZN(_1738_));
 AOI21_X1 _3919_ (.A(_1719_),
    .B1(_1727_),
    .B2(_1738_),
    .ZN(_0575_));
 NOR2_X1 _3920_ (.A1(prdata[30]),
    .A2(_1130_),
    .ZN(_1739_));
 AOI22_X1 _3921_ (.A1(\mem[18] [30]),
    .A2(net63),
    .B1(net36),
    .B2(\mem[23] [30]),
    .ZN(_1740_));
 AOI22_X1 _3922_ (.A1(\mem[11] [30]),
    .A2(net37),
    .B1(net20),
    .B2(\mem[8] [30]),
    .ZN(_1741_));
 AOI22_X1 _3923_ (.A1(\mem[12] [30]),
    .A2(net15),
    .B1(net5),
    .B2(\mem[9] [30]),
    .ZN(_1742_));
 AOI22_X1 _3924_ (.A1(\mem[14] [30]),
    .A2(net28),
    .B1(_1146_),
    .B2(\mem[25] [30]),
    .ZN(_1743_));
 AND4_X1 _3925_ (.A1(_1740_),
    .A2(_1741_),
    .A3(_1742_),
    .A4(_1743_),
    .ZN(_1744_));
 AOI222_X1 _3926_ (.A1(\mem[5] [30]),
    .A2(_1138_),
    .B1(_1147_),
    .B2(\mem[6] [30]),
    .C1(net24),
    .C2(\mem[1] [30]),
    .ZN(_1745_));
 AOI22_X1 _3927_ (.A1(\mem[26] [30]),
    .A2(_1096_),
    .B1(net44),
    .B2(\mem[3] [30]),
    .ZN(_1746_));
 AOI222_X1 _3928_ (.A1(\mem[15] [30]),
    .A2(net12),
    .B1(net53),
    .B2(\mem[20] [30]),
    .C1(_1128_),
    .C2(\mem[22] [30]),
    .ZN(_1747_));
 AOI222_X1 _3929_ (.A1(\mem[16] [30]),
    .A2(net9),
    .B1(_1105_),
    .B2(\mem[27] [30]),
    .C1(net51),
    .C2(\mem[2] [30]),
    .ZN(_1748_));
 NAND4_X1 _3930_ (.A1(_1745_),
    .A2(_1746_),
    .A3(_1747_),
    .A4(_1748_),
    .ZN(_1749_));
 AOI222_X1 _3931_ (.A1(\mem[0] [30]),
    .A2(net45),
    .B1(net41),
    .B2(\mem[4] [30]),
    .C1(net18),
    .C2(\mem[7] [30]),
    .ZN(_1750_));
 AOI221_X1 _3932_ (.A(net4),
    .B1(net47),
    .B2(\mem[30] [30]),
    .C1(\mem[31] [30]),
    .C2(net7),
    .ZN(_1751_));
 NAND2_X1 _3933_ (.A1(_1750_),
    .A2(_1751_),
    .ZN(_1752_));
 AOI22_X1 _3934_ (.A1(\mem[28] [30]),
    .A2(net61),
    .B1(net31),
    .B2(\mem[13] [30]),
    .ZN(_1753_));
 AOI22_X1 _3935_ (.A1(\mem[19] [30]),
    .A2(net59),
    .B1(_1135_),
    .B2(\mem[10] [30]),
    .ZN(_1754_));
 AOI22_X1 _3936_ (.A1(\mem[17] [30]),
    .A2(net70),
    .B1(_1123_),
    .B2(\mem[21] [30]),
    .ZN(_1755_));
 AOI22_X1 _3937_ (.A1(\mem[24] [30]),
    .A2(net56),
    .B1(net26),
    .B2(\mem[29] [30]),
    .ZN(_1756_));
 NAND4_X1 _3938_ (.A1(_1753_),
    .A2(_1754_),
    .A3(_1755_),
    .A4(_1756_),
    .ZN(_1757_));
 NOR3_X1 _3939_ (.A1(_1749_),
    .A2(_1752_),
    .A3(_1757_),
    .ZN(_1758_));
 AOI21_X1 _3940_ (.A(_1739_),
    .B1(_1744_),
    .B2(_1758_),
    .ZN(_0576_));
 NOR2_X1 _3941_ (.A1(prdata[31]),
    .A2(_1130_),
    .ZN(_1759_));
 AOI22_X1 _3942_ (.A1(\mem[5] [31]),
    .A2(_1138_),
    .B1(net17),
    .B2(\mem[7] [31]),
    .ZN(_1760_));
 AOI222_X1 _3943_ (.A1(\mem[26] [31]),
    .A2(_1096_),
    .B1(net51),
    .B2(\mem[2] [31]),
    .C1(net24),
    .C2(\mem[1] [31]),
    .ZN(_1761_));
 AOI221_X1 _3944_ (.A(net4),
    .B1(net36),
    .B2(\mem[23] [31]),
    .C1(_1123_),
    .C2(\mem[21] [31]),
    .ZN(_1762_));
 NAND2_X1 _3945_ (.A1(_1761_),
    .A2(_1762_),
    .ZN(_1763_));
 AOI22_X1 _3946_ (.A1(\mem[0] [31]),
    .A2(net45),
    .B1(_1147_),
    .B2(\mem[6] [31]),
    .ZN(_1764_));
 AOI22_X1 _3947_ (.A1(\mem[9] [31]),
    .A2(_1116_),
    .B1(net44),
    .B2(\mem[3] [31]),
    .ZN(_1765_));
 AOI22_X1 _3948_ (.A1(\mem[19] [31]),
    .A2(net60),
    .B1(_1146_),
    .B2(\mem[25] [31]),
    .ZN(_1766_));
 NAND4_X1 _3949_ (.A1(_1760_),
    .A2(_1764_),
    .A3(_1765_),
    .A4(_1766_),
    .ZN(_1767_));
 NOR2_X1 _3950_ (.A1(_1763_),
    .A2(_1767_),
    .ZN(_1768_));
 AOI222_X1 _3951_ (.A1(\mem[20] [31]),
    .A2(net55),
    .B1(_1135_),
    .B2(\mem[10] [31]),
    .C1(_1139_),
    .C2(\mem[11] [31]),
    .ZN(_1769_));
 AOI22_X1 _3952_ (.A1(\mem[16] [31]),
    .A2(net11),
    .B1(net66),
    .B2(\mem[27] [31]),
    .ZN(_1770_));
 AOI222_X2 _3953_ (.A1(\mem[12] [31]),
    .A2(_1077_),
    .B1(net68),
    .B2(\mem[17] [31]),
    .C1(net64),
    .C2(\mem[18] [31]),
    .ZN(_1771_));
 AOI222_X2 _3954_ (.A1(\mem[31] [31]),
    .A2(_1101_),
    .B1(net57),
    .B2(\mem[24] [31]),
    .C1(net21),
    .C2(\mem[8] [31]),
    .ZN(_1772_));
 NAND4_X1 _3955_ (.A1(_1769_),
    .A2(_1770_),
    .A3(_1771_),
    .A4(_1772_),
    .ZN(_1773_));
 AOI22_X1 _3956_ (.A1(\mem[4] [31]),
    .A2(net40),
    .B1(_1143_),
    .B2(\mem[29] [31]),
    .ZN(_1774_));
 AOI22_X1 _3957_ (.A1(\mem[22] [31]),
    .A2(_1128_),
    .B1(net27),
    .B2(\mem[14] [31]),
    .ZN(_1775_));
 AOI22_X1 _3958_ (.A1(\mem[28] [31]),
    .A2(net61),
    .B1(net47),
    .B2(\mem[30] [31]),
    .ZN(_1776_));
 AOI22_X1 _3959_ (.A1(\mem[15] [31]),
    .A2(net13),
    .B1(net32),
    .B2(\mem[13] [31]),
    .ZN(_1777_));
 NAND4_X1 _3960_ (.A1(_1774_),
    .A2(_1775_),
    .A3(_1776_),
    .A4(_1777_),
    .ZN(_1778_));
 NOR2_X1 _3961_ (.A1(_1773_),
    .A2(_1778_),
    .ZN(_1779_));
 AOI21_X1 _3962_ (.A(_1759_),
    .B1(_1768_),
    .B2(_1779_),
    .ZN(_0577_));
 NAND2_X4 _3963_ (.A1(net2),
    .A2(net23),
    .ZN(_1780_));
 MUX2_X1 _3964_ (.A(pwdata[0]),
    .B(\mem[1] [0]),
    .S(_1780_),
    .Z(_0578_));
 MUX2_X1 _3965_ (.A(pwdata[1]),
    .B(\mem[1] [1]),
    .S(_1780_),
    .Z(_0579_));
 MUX2_X1 _3966_ (.A(pwdata[2]),
    .B(\mem[1] [2]),
    .S(_1780_),
    .Z(_0580_));
 MUX2_X1 _3967_ (.A(pwdata[3]),
    .B(\mem[1] [3]),
    .S(_1780_),
    .Z(_0581_));
 MUX2_X1 _3968_ (.A(pwdata[4]),
    .B(\mem[1] [4]),
    .S(_1780_),
    .Z(_0582_));
 MUX2_X1 _3969_ (.A(pwdata[5]),
    .B(\mem[1] [5]),
    .S(_1780_),
    .Z(_0583_));
 MUX2_X1 _3970_ (.A(pwdata[6]),
    .B(\mem[1] [6]),
    .S(_1780_),
    .Z(_0584_));
 MUX2_X1 _3971_ (.A(pwdata[7]),
    .B(\mem[1] [7]),
    .S(_1780_),
    .Z(_0585_));
 MUX2_X1 _3972_ (.A(pwdata[8]),
    .B(\mem[1] [8]),
    .S(_1780_),
    .Z(_0586_));
 MUX2_X1 _3973_ (.A(pwdata[9]),
    .B(\mem[1] [9]),
    .S(_1780_),
    .Z(_0587_));
 MUX2_X1 _3974_ (.A(pwdata[10]),
    .B(\mem[1] [10]),
    .S(_1780_),
    .Z(_0588_));
 MUX2_X1 _3975_ (.A(pwdata[11]),
    .B(\mem[1] [11]),
    .S(_1780_),
    .Z(_0589_));
 MUX2_X1 _3976_ (.A(pwdata[12]),
    .B(\mem[1] [12]),
    .S(_1780_),
    .Z(_0590_));
 MUX2_X1 _3977_ (.A(pwdata[13]),
    .B(\mem[1] [13]),
    .S(_1780_),
    .Z(_0591_));
 MUX2_X1 _3978_ (.A(pwdata[14]),
    .B(\mem[1] [14]),
    .S(_1780_),
    .Z(_0592_));
 MUX2_X1 _3979_ (.A(pwdata[15]),
    .B(\mem[1] [15]),
    .S(_1780_),
    .Z(_0593_));
 MUX2_X1 _3980_ (.A(pwdata[16]),
    .B(\mem[1] [16]),
    .S(_1780_),
    .Z(_0594_));
 MUX2_X1 _3981_ (.A(pwdata[17]),
    .B(\mem[1] [17]),
    .S(_1780_),
    .Z(_0595_));
 MUX2_X1 _3982_ (.A(pwdata[18]),
    .B(\mem[1] [18]),
    .S(_1780_),
    .Z(_0596_));
 MUX2_X1 _3983_ (.A(pwdata[19]),
    .B(\mem[1] [19]),
    .S(_1780_),
    .Z(_0597_));
 MUX2_X1 _3984_ (.A(pwdata[20]),
    .B(\mem[1] [20]),
    .S(_1780_),
    .Z(_0598_));
 MUX2_X1 _3985_ (.A(pwdata[21]),
    .B(\mem[1] [21]),
    .S(_1780_),
    .Z(_0599_));
 MUX2_X1 _3986_ (.A(pwdata[22]),
    .B(\mem[1] [22]),
    .S(_1780_),
    .Z(_0600_));
 MUX2_X1 _3987_ (.A(pwdata[23]),
    .B(\mem[1] [23]),
    .S(_1780_),
    .Z(_0601_));
 MUX2_X1 _3988_ (.A(pwdata[24]),
    .B(\mem[1] [24]),
    .S(_1780_),
    .Z(_0602_));
 MUX2_X1 _3989_ (.A(pwdata[25]),
    .B(\mem[1] [25]),
    .S(_1780_),
    .Z(_0603_));
 MUX2_X1 _3990_ (.A(pwdata[26]),
    .B(\mem[1] [26]),
    .S(_1780_),
    .Z(_0604_));
 MUX2_X1 _3991_ (.A(pwdata[27]),
    .B(\mem[1] [27]),
    .S(_1780_),
    .Z(_0605_));
 MUX2_X1 _3992_ (.A(pwdata[28]),
    .B(\mem[1] [28]),
    .S(_1780_),
    .Z(_0606_));
 MUX2_X1 _3993_ (.A(pwdata[29]),
    .B(\mem[1] [29]),
    .S(_1780_),
    .Z(_0607_));
 MUX2_X1 _3994_ (.A(pwdata[30]),
    .B(\mem[1] [30]),
    .S(_1780_),
    .Z(_0608_));
 MUX2_X1 _3995_ (.A(pwdata[31]),
    .B(\mem[1] [31]),
    .S(_1780_),
    .Z(_0609_));
 NAND2_X4 _3996_ (.A1(net2),
    .A2(net35),
    .ZN(_1781_));
 MUX2_X1 _3997_ (.A(pwdata[0]),
    .B(\mem[23] [0]),
    .S(_1781_),
    .Z(_0610_));
 MUX2_X1 _3998_ (.A(pwdata[1]),
    .B(\mem[23] [1]),
    .S(_1781_),
    .Z(_0611_));
 MUX2_X1 _3999_ (.A(pwdata[2]),
    .B(\mem[23] [2]),
    .S(_1781_),
    .Z(_0612_));
 MUX2_X1 _4000_ (.A(pwdata[3]),
    .B(\mem[23] [3]),
    .S(_1781_),
    .Z(_0613_));
 MUX2_X1 _4001_ (.A(pwdata[4]),
    .B(\mem[23] [4]),
    .S(_1781_),
    .Z(_0614_));
 MUX2_X1 _4002_ (.A(pwdata[5]),
    .B(\mem[23] [5]),
    .S(_1781_),
    .Z(_0615_));
 MUX2_X1 _4003_ (.A(pwdata[6]),
    .B(\mem[23] [6]),
    .S(_1781_),
    .Z(_0616_));
 MUX2_X1 _4004_ (.A(pwdata[7]),
    .B(\mem[23] [7]),
    .S(_1781_),
    .Z(_0617_));
 MUX2_X1 _4005_ (.A(pwdata[8]),
    .B(\mem[23] [8]),
    .S(_1781_),
    .Z(_0618_));
 MUX2_X1 _4006_ (.A(pwdata[9]),
    .B(\mem[23] [9]),
    .S(_1781_),
    .Z(_0619_));
 MUX2_X1 _4007_ (.A(pwdata[10]),
    .B(\mem[23] [10]),
    .S(_1781_),
    .Z(_0620_));
 MUX2_X1 _4008_ (.A(pwdata[11]),
    .B(\mem[23] [11]),
    .S(_1781_),
    .Z(_0621_));
 MUX2_X1 _4009_ (.A(pwdata[12]),
    .B(\mem[23] [12]),
    .S(_1781_),
    .Z(_0622_));
 MUX2_X1 _4010_ (.A(pwdata[13]),
    .B(\mem[23] [13]),
    .S(_1781_),
    .Z(_0623_));
 MUX2_X1 _4011_ (.A(pwdata[14]),
    .B(\mem[23] [14]),
    .S(_1781_),
    .Z(_0624_));
 MUX2_X1 _4012_ (.A(pwdata[15]),
    .B(\mem[23] [15]),
    .S(_1781_),
    .Z(_0625_));
 MUX2_X1 _4013_ (.A(pwdata[16]),
    .B(\mem[23] [16]),
    .S(_1781_),
    .Z(_0626_));
 MUX2_X1 _4014_ (.A(pwdata[17]),
    .B(\mem[23] [17]),
    .S(_1781_),
    .Z(_0627_));
 MUX2_X1 _4015_ (.A(pwdata[18]),
    .B(\mem[23] [18]),
    .S(_1781_),
    .Z(_0628_));
 MUX2_X1 _4016_ (.A(pwdata[19]),
    .B(\mem[23] [19]),
    .S(_1781_),
    .Z(_0629_));
 MUX2_X1 _4017_ (.A(pwdata[20]),
    .B(\mem[23] [20]),
    .S(_1781_),
    .Z(_0630_));
 MUX2_X1 _4018_ (.A(pwdata[21]),
    .B(\mem[23] [21]),
    .S(_1781_),
    .Z(_0631_));
 MUX2_X1 _4019_ (.A(pwdata[22]),
    .B(\mem[23] [22]),
    .S(_1781_),
    .Z(_0632_));
 MUX2_X1 _4020_ (.A(pwdata[23]),
    .B(\mem[23] [23]),
    .S(_1781_),
    .Z(_0633_));
 MUX2_X1 _4021_ (.A(pwdata[24]),
    .B(\mem[23] [24]),
    .S(_1781_),
    .Z(_0634_));
 MUX2_X1 _4022_ (.A(pwdata[25]),
    .B(\mem[23] [25]),
    .S(_1781_),
    .Z(_0635_));
 MUX2_X1 _4023_ (.A(pwdata[26]),
    .B(\mem[23] [26]),
    .S(_1781_),
    .Z(_0636_));
 MUX2_X1 _4024_ (.A(pwdata[27]),
    .B(\mem[23] [27]),
    .S(_1781_),
    .Z(_0637_));
 MUX2_X1 _4025_ (.A(pwdata[28]),
    .B(\mem[23] [28]),
    .S(_1781_),
    .Z(_0638_));
 MUX2_X1 _4026_ (.A(pwdata[29]),
    .B(\mem[23] [29]),
    .S(_1781_),
    .Z(_0639_));
 MUX2_X1 _4027_ (.A(pwdata[30]),
    .B(\mem[23] [30]),
    .S(_1781_),
    .Z(_0640_));
 MUX2_X1 _4028_ (.A(pwdata[31]),
    .B(\mem[23] [31]),
    .S(_1781_),
    .Z(_0641_));
 NAND2_X4 _4029_ (.A1(net2),
    .A2(_1146_),
    .ZN(_1782_));
 MUX2_X1 _4030_ (.A(pwdata[0]),
    .B(\mem[25] [0]),
    .S(_1782_),
    .Z(_0642_));
 MUX2_X1 _4031_ (.A(pwdata[1]),
    .B(\mem[25] [1]),
    .S(_1782_),
    .Z(_0643_));
 MUX2_X1 _4032_ (.A(pwdata[2]),
    .B(\mem[25] [2]),
    .S(_1782_),
    .Z(_0644_));
 MUX2_X1 _4033_ (.A(pwdata[3]),
    .B(\mem[25] [3]),
    .S(_1782_),
    .Z(_0645_));
 MUX2_X1 _4034_ (.A(pwdata[4]),
    .B(\mem[25] [4]),
    .S(_1782_),
    .Z(_0646_));
 MUX2_X1 _4035_ (.A(pwdata[5]),
    .B(\mem[25] [5]),
    .S(_1782_),
    .Z(_0647_));
 MUX2_X1 _4036_ (.A(pwdata[6]),
    .B(\mem[25] [6]),
    .S(_1782_),
    .Z(_0648_));
 MUX2_X1 _4037_ (.A(pwdata[7]),
    .B(\mem[25] [7]),
    .S(_1782_),
    .Z(_0649_));
 MUX2_X1 _4038_ (.A(pwdata[8]),
    .B(\mem[25] [8]),
    .S(_1782_),
    .Z(_0650_));
 MUX2_X1 _4039_ (.A(pwdata[9]),
    .B(\mem[25] [9]),
    .S(_1782_),
    .Z(_0651_));
 MUX2_X1 _4040_ (.A(pwdata[10]),
    .B(\mem[25] [10]),
    .S(_1782_),
    .Z(_0652_));
 MUX2_X1 _4041_ (.A(pwdata[11]),
    .B(\mem[25] [11]),
    .S(_1782_),
    .Z(_0653_));
 MUX2_X1 _4042_ (.A(pwdata[12]),
    .B(\mem[25] [12]),
    .S(_1782_),
    .Z(_0654_));
 MUX2_X1 _4043_ (.A(pwdata[13]),
    .B(\mem[25] [13]),
    .S(_1782_),
    .Z(_0655_));
 MUX2_X1 _4044_ (.A(pwdata[14]),
    .B(\mem[25] [14]),
    .S(_1782_),
    .Z(_0656_));
 MUX2_X1 _4045_ (.A(pwdata[15]),
    .B(\mem[25] [15]),
    .S(_1782_),
    .Z(_0657_));
 MUX2_X1 _4046_ (.A(pwdata[16]),
    .B(\mem[25] [16]),
    .S(_1782_),
    .Z(_0658_));
 MUX2_X1 _4047_ (.A(pwdata[17]),
    .B(\mem[25] [17]),
    .S(_1782_),
    .Z(_0659_));
 MUX2_X1 _4048_ (.A(pwdata[18]),
    .B(\mem[25] [18]),
    .S(_1782_),
    .Z(_0660_));
 MUX2_X1 _4049_ (.A(pwdata[19]),
    .B(\mem[25] [19]),
    .S(_1782_),
    .Z(_0661_));
 MUX2_X1 _4050_ (.A(pwdata[20]),
    .B(\mem[25] [20]),
    .S(_1782_),
    .Z(_0662_));
 MUX2_X1 _4051_ (.A(pwdata[21]),
    .B(\mem[25] [21]),
    .S(_1782_),
    .Z(_0663_));
 MUX2_X1 _4052_ (.A(pwdata[22]),
    .B(\mem[25] [22]),
    .S(_1782_),
    .Z(_0664_));
 MUX2_X1 _4053_ (.A(pwdata[23]),
    .B(\mem[25] [23]),
    .S(_1782_),
    .Z(_0665_));
 MUX2_X1 _4054_ (.A(pwdata[24]),
    .B(\mem[25] [24]),
    .S(_1782_),
    .Z(_0666_));
 MUX2_X1 _4055_ (.A(pwdata[25]),
    .B(\mem[25] [25]),
    .S(_1782_),
    .Z(_0667_));
 MUX2_X1 _4056_ (.A(pwdata[26]),
    .B(\mem[25] [26]),
    .S(_1782_),
    .Z(_0668_));
 MUX2_X1 _4057_ (.A(pwdata[27]),
    .B(\mem[25] [27]),
    .S(_1782_),
    .Z(_0669_));
 MUX2_X1 _4058_ (.A(pwdata[28]),
    .B(\mem[25] [28]),
    .S(_1782_),
    .Z(_0670_));
 MUX2_X1 _4059_ (.A(pwdata[29]),
    .B(\mem[25] [29]),
    .S(_1782_),
    .Z(_0671_));
 MUX2_X1 _4060_ (.A(pwdata[30]),
    .B(\mem[25] [30]),
    .S(_1782_),
    .Z(_0672_));
 MUX2_X1 _4061_ (.A(pwdata[31]),
    .B(\mem[25] [31]),
    .S(_1782_),
    .Z(_0673_));
 NAND2_X4 _4062_ (.A1(net2),
    .A2(net16),
    .ZN(_1783_));
 MUX2_X1 _4063_ (.A(pwdata[0]),
    .B(\mem[7] [0]),
    .S(_1783_),
    .Z(_0674_));
 MUX2_X1 _4064_ (.A(pwdata[1]),
    .B(\mem[7] [1]),
    .S(_1783_),
    .Z(_0675_));
 MUX2_X1 _4065_ (.A(pwdata[2]),
    .B(\mem[7] [2]),
    .S(_1783_),
    .Z(_0676_));
 MUX2_X1 _4066_ (.A(pwdata[3]),
    .B(\mem[7] [3]),
    .S(_1783_),
    .Z(_0677_));
 MUX2_X1 _4067_ (.A(pwdata[4]),
    .B(\mem[7] [4]),
    .S(_1783_),
    .Z(_0678_));
 MUX2_X1 _4068_ (.A(pwdata[5]),
    .B(\mem[7] [5]),
    .S(_1783_),
    .Z(_0679_));
 MUX2_X1 _4069_ (.A(pwdata[6]),
    .B(\mem[7] [6]),
    .S(_1783_),
    .Z(_0680_));
 MUX2_X1 _4070_ (.A(pwdata[7]),
    .B(\mem[7] [7]),
    .S(_1783_),
    .Z(_0681_));
 MUX2_X1 _4071_ (.A(pwdata[8]),
    .B(\mem[7] [8]),
    .S(_1783_),
    .Z(_0682_));
 MUX2_X1 _4072_ (.A(pwdata[9]),
    .B(\mem[7] [9]),
    .S(_1783_),
    .Z(_0683_));
 MUX2_X1 _4073_ (.A(pwdata[10]),
    .B(\mem[7] [10]),
    .S(_1783_),
    .Z(_0684_));
 MUX2_X1 _4074_ (.A(pwdata[11]),
    .B(\mem[7] [11]),
    .S(_1783_),
    .Z(_0685_));
 MUX2_X1 _4075_ (.A(pwdata[12]),
    .B(\mem[7] [12]),
    .S(_1783_),
    .Z(_0686_));
 MUX2_X1 _4076_ (.A(pwdata[13]),
    .B(\mem[7] [13]),
    .S(_1783_),
    .Z(_0687_));
 MUX2_X1 _4077_ (.A(pwdata[14]),
    .B(\mem[7] [14]),
    .S(_1783_),
    .Z(_0688_));
 MUX2_X1 _4078_ (.A(pwdata[15]),
    .B(\mem[7] [15]),
    .S(_1783_),
    .Z(_0689_));
 MUX2_X1 _4079_ (.A(pwdata[16]),
    .B(\mem[7] [16]),
    .S(_1783_),
    .Z(_0690_));
 MUX2_X1 _4080_ (.A(pwdata[17]),
    .B(\mem[7] [17]),
    .S(_1783_),
    .Z(_0691_));
 MUX2_X1 _4081_ (.A(pwdata[18]),
    .B(\mem[7] [18]),
    .S(_1783_),
    .Z(_0692_));
 MUX2_X1 _4082_ (.A(pwdata[19]),
    .B(\mem[7] [19]),
    .S(_1783_),
    .Z(_0693_));
 MUX2_X1 _4083_ (.A(pwdata[20]),
    .B(\mem[7] [20]),
    .S(_1783_),
    .Z(_0694_));
 MUX2_X1 _4084_ (.A(pwdata[21]),
    .B(\mem[7] [21]),
    .S(_1783_),
    .Z(_0695_));
 MUX2_X1 _4085_ (.A(pwdata[22]),
    .B(\mem[7] [22]),
    .S(_1783_),
    .Z(_0696_));
 MUX2_X1 _4086_ (.A(pwdata[23]),
    .B(\mem[7] [23]),
    .S(_1783_),
    .Z(_0697_));
 MUX2_X1 _4087_ (.A(pwdata[24]),
    .B(\mem[7] [24]),
    .S(_1783_),
    .Z(_0698_));
 MUX2_X1 _4088_ (.A(pwdata[25]),
    .B(\mem[7] [25]),
    .S(_1783_),
    .Z(_0699_));
 MUX2_X1 _4089_ (.A(pwdata[26]),
    .B(\mem[7] [26]),
    .S(_1783_),
    .Z(_0700_));
 MUX2_X1 _4090_ (.A(pwdata[27]),
    .B(\mem[7] [27]),
    .S(_1783_),
    .Z(_0701_));
 MUX2_X1 _4091_ (.A(pwdata[28]),
    .B(\mem[7] [28]),
    .S(_1783_),
    .Z(_0702_));
 MUX2_X1 _4092_ (.A(pwdata[29]),
    .B(\mem[7] [29]),
    .S(_1783_),
    .Z(_0703_));
 MUX2_X1 _4093_ (.A(pwdata[30]),
    .B(\mem[7] [30]),
    .S(_1783_),
    .Z(_0704_));
 MUX2_X1 _4094_ (.A(pwdata[31]),
    .B(\mem[7] [31]),
    .S(_1783_),
    .Z(_0705_));
 NAND2_X4 _4095_ (.A1(net2),
    .A2(_1135_),
    .ZN(_1784_));
 MUX2_X1 _4096_ (.A(pwdata[0]),
    .B(\mem[10] [0]),
    .S(_1784_),
    .Z(_0706_));
 MUX2_X1 _4097_ (.A(pwdata[1]),
    .B(\mem[10] [1]),
    .S(_1784_),
    .Z(_0707_));
 MUX2_X1 _4098_ (.A(pwdata[2]),
    .B(\mem[10] [2]),
    .S(_1784_),
    .Z(_0708_));
 MUX2_X1 _4099_ (.A(pwdata[3]),
    .B(\mem[10] [3]),
    .S(_1784_),
    .Z(_0709_));
 MUX2_X1 _4100_ (.A(pwdata[4]),
    .B(\mem[10] [4]),
    .S(_1784_),
    .Z(_0710_));
 MUX2_X1 _4101_ (.A(pwdata[5]),
    .B(\mem[10] [5]),
    .S(_1784_),
    .Z(_0711_));
 MUX2_X1 _4102_ (.A(pwdata[6]),
    .B(\mem[10] [6]),
    .S(_1784_),
    .Z(_0712_));
 MUX2_X1 _4103_ (.A(pwdata[7]),
    .B(\mem[10] [7]),
    .S(_1784_),
    .Z(_0713_));
 MUX2_X1 _4104_ (.A(pwdata[8]),
    .B(\mem[10] [8]),
    .S(_1784_),
    .Z(_0714_));
 MUX2_X1 _4105_ (.A(pwdata[9]),
    .B(\mem[10] [9]),
    .S(_1784_),
    .Z(_0715_));
 MUX2_X1 _4106_ (.A(pwdata[10]),
    .B(\mem[10] [10]),
    .S(_1784_),
    .Z(_0716_));
 MUX2_X1 _4107_ (.A(pwdata[11]),
    .B(\mem[10] [11]),
    .S(_1784_),
    .Z(_0717_));
 MUX2_X1 _4108_ (.A(pwdata[12]),
    .B(\mem[10] [12]),
    .S(_1784_),
    .Z(_0718_));
 MUX2_X1 _4109_ (.A(pwdata[13]),
    .B(\mem[10] [13]),
    .S(_1784_),
    .Z(_0719_));
 MUX2_X1 _4110_ (.A(pwdata[14]),
    .B(\mem[10] [14]),
    .S(_1784_),
    .Z(_0720_));
 MUX2_X1 _4111_ (.A(pwdata[15]),
    .B(\mem[10] [15]),
    .S(_1784_),
    .Z(_0721_));
 MUX2_X1 _4112_ (.A(pwdata[16]),
    .B(\mem[10] [16]),
    .S(_1784_),
    .Z(_0722_));
 MUX2_X1 _4113_ (.A(pwdata[17]),
    .B(\mem[10] [17]),
    .S(_1784_),
    .Z(_0723_));
 MUX2_X1 _4114_ (.A(pwdata[18]),
    .B(\mem[10] [18]),
    .S(_1784_),
    .Z(_0724_));
 MUX2_X1 _4115_ (.A(pwdata[19]),
    .B(\mem[10] [19]),
    .S(_1784_),
    .Z(_0725_));
 MUX2_X1 _4116_ (.A(pwdata[20]),
    .B(\mem[10] [20]),
    .S(_1784_),
    .Z(_0726_));
 MUX2_X1 _4117_ (.A(pwdata[21]),
    .B(\mem[10] [21]),
    .S(_1784_),
    .Z(_0727_));
 MUX2_X1 _4118_ (.A(pwdata[22]),
    .B(\mem[10] [22]),
    .S(_1784_),
    .Z(_0728_));
 MUX2_X1 _4119_ (.A(pwdata[23]),
    .B(\mem[10] [23]),
    .S(_1784_),
    .Z(_0729_));
 MUX2_X1 _4120_ (.A(pwdata[24]),
    .B(\mem[10] [24]),
    .S(_1784_),
    .Z(_0730_));
 MUX2_X1 _4121_ (.A(pwdata[25]),
    .B(\mem[10] [25]),
    .S(_1784_),
    .Z(_0731_));
 MUX2_X1 _4122_ (.A(pwdata[26]),
    .B(\mem[10] [26]),
    .S(_1784_),
    .Z(_0732_));
 MUX2_X1 _4123_ (.A(pwdata[27]),
    .B(\mem[10] [27]),
    .S(_1784_),
    .Z(_0733_));
 MUX2_X1 _4124_ (.A(pwdata[28]),
    .B(\mem[10] [28]),
    .S(_1784_),
    .Z(_0734_));
 MUX2_X1 _4125_ (.A(pwdata[29]),
    .B(\mem[10] [29]),
    .S(_1784_),
    .Z(_0735_));
 MUX2_X1 _4126_ (.A(pwdata[30]),
    .B(\mem[10] [30]),
    .S(_1784_),
    .Z(_0736_));
 MUX2_X1 _4127_ (.A(pwdata[31]),
    .B(\mem[10] [31]),
    .S(_1784_),
    .Z(_0737_));
 NAND2_X4 _4128_ (.A1(net2),
    .A2(net26),
    .ZN(_1785_));
 MUX2_X1 _4129_ (.A(pwdata[0]),
    .B(\mem[29] [0]),
    .S(_1785_),
    .Z(_0738_));
 MUX2_X1 _4130_ (.A(pwdata[1]),
    .B(\mem[29] [1]),
    .S(_1785_),
    .Z(_0739_));
 MUX2_X1 _4131_ (.A(pwdata[2]),
    .B(\mem[29] [2]),
    .S(_1785_),
    .Z(_0740_));
 MUX2_X1 _4132_ (.A(pwdata[3]),
    .B(\mem[29] [3]),
    .S(_1785_),
    .Z(_0741_));
 MUX2_X1 _4133_ (.A(pwdata[4]),
    .B(\mem[29] [4]),
    .S(_1785_),
    .Z(_0742_));
 MUX2_X1 _4134_ (.A(pwdata[5]),
    .B(\mem[29] [5]),
    .S(_1785_),
    .Z(_0743_));
 MUX2_X1 _4135_ (.A(pwdata[6]),
    .B(\mem[29] [6]),
    .S(_1785_),
    .Z(_0744_));
 MUX2_X1 _4136_ (.A(pwdata[7]),
    .B(\mem[29] [7]),
    .S(_1785_),
    .Z(_0745_));
 MUX2_X1 _4137_ (.A(pwdata[8]),
    .B(\mem[29] [8]),
    .S(_1785_),
    .Z(_0746_));
 MUX2_X1 _4138_ (.A(pwdata[9]),
    .B(\mem[29] [9]),
    .S(_1785_),
    .Z(_0747_));
 MUX2_X1 _4139_ (.A(pwdata[10]),
    .B(\mem[29] [10]),
    .S(_1785_),
    .Z(_0748_));
 MUX2_X1 _4140_ (.A(pwdata[11]),
    .B(\mem[29] [11]),
    .S(_1785_),
    .Z(_0749_));
 MUX2_X1 _4141_ (.A(pwdata[12]),
    .B(\mem[29] [12]),
    .S(_1785_),
    .Z(_0750_));
 MUX2_X1 _4142_ (.A(pwdata[13]),
    .B(\mem[29] [13]),
    .S(_1785_),
    .Z(_0751_));
 MUX2_X1 _4143_ (.A(pwdata[14]),
    .B(\mem[29] [14]),
    .S(_1785_),
    .Z(_0752_));
 MUX2_X1 _4144_ (.A(pwdata[15]),
    .B(\mem[29] [15]),
    .S(_1785_),
    .Z(_0753_));
 MUX2_X1 _4145_ (.A(pwdata[16]),
    .B(\mem[29] [16]),
    .S(_1785_),
    .Z(_0754_));
 MUX2_X1 _4146_ (.A(pwdata[17]),
    .B(\mem[29] [17]),
    .S(_1785_),
    .Z(_0755_));
 MUX2_X1 _4147_ (.A(pwdata[18]),
    .B(\mem[29] [18]),
    .S(_1785_),
    .Z(_0756_));
 MUX2_X1 _4148_ (.A(pwdata[19]),
    .B(\mem[29] [19]),
    .S(_1785_),
    .Z(_0757_));
 MUX2_X1 _4149_ (.A(pwdata[20]),
    .B(\mem[29] [20]),
    .S(_1785_),
    .Z(_0758_));
 MUX2_X1 _4150_ (.A(pwdata[21]),
    .B(\mem[29] [21]),
    .S(_1785_),
    .Z(_0759_));
 MUX2_X1 _4151_ (.A(pwdata[22]),
    .B(\mem[29] [22]),
    .S(_1785_),
    .Z(_0760_));
 MUX2_X1 _4152_ (.A(pwdata[23]),
    .B(\mem[29] [23]),
    .S(_1785_),
    .Z(_0761_));
 MUX2_X1 _4153_ (.A(pwdata[24]),
    .B(\mem[29] [24]),
    .S(_1785_),
    .Z(_0762_));
 MUX2_X1 _4154_ (.A(pwdata[25]),
    .B(\mem[29] [25]),
    .S(_1785_),
    .Z(_0763_));
 MUX2_X1 _4155_ (.A(pwdata[26]),
    .B(\mem[29] [26]),
    .S(_1785_),
    .Z(_0764_));
 MUX2_X1 _4156_ (.A(pwdata[27]),
    .B(\mem[29] [27]),
    .S(_1785_),
    .Z(_0765_));
 MUX2_X1 _4157_ (.A(pwdata[28]),
    .B(\mem[29] [28]),
    .S(_1785_),
    .Z(_0766_));
 MUX2_X1 _4158_ (.A(pwdata[29]),
    .B(\mem[29] [29]),
    .S(_1785_),
    .Z(_0767_));
 MUX2_X1 _4159_ (.A(pwdata[30]),
    .B(\mem[29] [30]),
    .S(_1785_),
    .Z(_0768_));
 MUX2_X1 _4160_ (.A(pwdata[31]),
    .B(\mem[29] [31]),
    .S(_1785_),
    .Z(_0769_));
 AOI21_X1 _4161_ (.A(_1089_),
    .B1(_1083_),
    .B2(_1068_),
    .ZN(_0770_));
 NAND2_X4 _4162_ (.A1(_1090_),
    .A2(net43),
    .ZN(_1786_));
 MUX2_X1 _4163_ (.A(pwdata[0]),
    .B(\mem[3] [0]),
    .S(_1786_),
    .Z(_0771_));
 MUX2_X1 _4164_ (.A(pwdata[1]),
    .B(\mem[3] [1]),
    .S(_1786_),
    .Z(_0772_));
 MUX2_X1 _4165_ (.A(pwdata[2]),
    .B(\mem[3] [2]),
    .S(_1786_),
    .Z(_0773_));
 MUX2_X1 _4166_ (.A(pwdata[3]),
    .B(\mem[3] [3]),
    .S(_1786_),
    .Z(_0774_));
 MUX2_X1 _4167_ (.A(pwdata[4]),
    .B(\mem[3] [4]),
    .S(_1786_),
    .Z(_0775_));
 MUX2_X1 _4168_ (.A(pwdata[5]),
    .B(\mem[3] [5]),
    .S(_1786_),
    .Z(_0776_));
 MUX2_X1 _4169_ (.A(pwdata[6]),
    .B(\mem[3] [6]),
    .S(_1786_),
    .Z(_0777_));
 MUX2_X1 _4170_ (.A(pwdata[7]),
    .B(\mem[3] [7]),
    .S(_1786_),
    .Z(_0778_));
 MUX2_X1 _4171_ (.A(pwdata[8]),
    .B(\mem[3] [8]),
    .S(_1786_),
    .Z(_0779_));
 MUX2_X1 _4172_ (.A(pwdata[9]),
    .B(\mem[3] [9]),
    .S(_1786_),
    .Z(_0780_));
 MUX2_X1 _4173_ (.A(pwdata[10]),
    .B(\mem[3] [10]),
    .S(_1786_),
    .Z(_0781_));
 MUX2_X1 _4174_ (.A(pwdata[11]),
    .B(\mem[3] [11]),
    .S(_1786_),
    .Z(_0782_));
 MUX2_X1 _4175_ (.A(pwdata[12]),
    .B(\mem[3] [12]),
    .S(_1786_),
    .Z(_0783_));
 MUX2_X1 _4176_ (.A(pwdata[13]),
    .B(\mem[3] [13]),
    .S(_1786_),
    .Z(_0784_));
 MUX2_X1 _4177_ (.A(pwdata[14]),
    .B(\mem[3] [14]),
    .S(_1786_),
    .Z(_0785_));
 MUX2_X1 _4178_ (.A(pwdata[15]),
    .B(\mem[3] [15]),
    .S(_1786_),
    .Z(_0786_));
 MUX2_X1 _4179_ (.A(pwdata[16]),
    .B(\mem[3] [16]),
    .S(_1786_),
    .Z(_0787_));
 MUX2_X1 _4180_ (.A(pwdata[17]),
    .B(\mem[3] [17]),
    .S(_1786_),
    .Z(_0788_));
 MUX2_X1 _4181_ (.A(pwdata[18]),
    .B(\mem[3] [18]),
    .S(_1786_),
    .Z(_0789_));
 MUX2_X1 _4182_ (.A(pwdata[19]),
    .B(\mem[3] [19]),
    .S(_1786_),
    .Z(_0790_));
 MUX2_X1 _4183_ (.A(pwdata[20]),
    .B(\mem[3] [20]),
    .S(_1786_),
    .Z(_0791_));
 MUX2_X1 _4184_ (.A(pwdata[21]),
    .B(\mem[3] [21]),
    .S(_1786_),
    .Z(_0792_));
 MUX2_X1 _4185_ (.A(pwdata[22]),
    .B(\mem[3] [22]),
    .S(_1786_),
    .Z(_0793_));
 MUX2_X1 _4186_ (.A(pwdata[23]),
    .B(\mem[3] [23]),
    .S(_1786_),
    .Z(_0794_));
 MUX2_X1 _4187_ (.A(pwdata[24]),
    .B(\mem[3] [24]),
    .S(_1786_),
    .Z(_0795_));
 MUX2_X1 _4188_ (.A(pwdata[25]),
    .B(\mem[3] [25]),
    .S(_1786_),
    .Z(_0796_));
 MUX2_X1 _4189_ (.A(pwdata[26]),
    .B(\mem[3] [26]),
    .S(_1786_),
    .Z(_0797_));
 MUX2_X1 _4190_ (.A(pwdata[27]),
    .B(\mem[3] [27]),
    .S(_1786_),
    .Z(_0798_));
 MUX2_X1 _4191_ (.A(pwdata[28]),
    .B(\mem[3] [28]),
    .S(_1786_),
    .Z(_0799_));
 MUX2_X1 _4192_ (.A(pwdata[29]),
    .B(\mem[3] [29]),
    .S(_1786_),
    .Z(_0800_));
 MUX2_X1 _4193_ (.A(pwdata[30]),
    .B(\mem[3] [30]),
    .S(_1786_),
    .Z(_0801_));
 MUX2_X1 _4194_ (.A(pwdata[31]),
    .B(\mem[3] [31]),
    .S(_1786_),
    .Z(_0802_));
 NAND2_X4 _4195_ (.A1(net2),
    .A2(net19),
    .ZN(_1787_));
 MUX2_X1 _4196_ (.A(pwdata[0]),
    .B(\mem[8] [0]),
    .S(_1787_),
    .Z(_0803_));
 MUX2_X1 _4197_ (.A(pwdata[1]),
    .B(\mem[8] [1]),
    .S(_1787_),
    .Z(_0804_));
 MUX2_X1 _4198_ (.A(pwdata[2]),
    .B(\mem[8] [2]),
    .S(_1787_),
    .Z(_0805_));
 MUX2_X1 _4199_ (.A(pwdata[3]),
    .B(\mem[8] [3]),
    .S(_1787_),
    .Z(_0806_));
 MUX2_X1 _4200_ (.A(pwdata[4]),
    .B(\mem[8] [4]),
    .S(_1787_),
    .Z(_0807_));
 MUX2_X1 _4201_ (.A(pwdata[5]),
    .B(\mem[8] [5]),
    .S(_1787_),
    .Z(_0808_));
 MUX2_X1 _4202_ (.A(pwdata[6]),
    .B(\mem[8] [6]),
    .S(_1787_),
    .Z(_0809_));
 MUX2_X1 _4203_ (.A(pwdata[7]),
    .B(\mem[8] [7]),
    .S(_1787_),
    .Z(_0810_));
 MUX2_X1 _4204_ (.A(pwdata[8]),
    .B(\mem[8] [8]),
    .S(_1787_),
    .Z(_0811_));
 MUX2_X1 _4205_ (.A(pwdata[9]),
    .B(\mem[8] [9]),
    .S(_1787_),
    .Z(_0812_));
 MUX2_X1 _4206_ (.A(pwdata[10]),
    .B(\mem[8] [10]),
    .S(_1787_),
    .Z(_0813_));
 MUX2_X1 _4207_ (.A(pwdata[11]),
    .B(\mem[8] [11]),
    .S(_1787_),
    .Z(_0814_));
 MUX2_X1 _4208_ (.A(pwdata[12]),
    .B(\mem[8] [12]),
    .S(_1787_),
    .Z(_0815_));
 MUX2_X1 _4209_ (.A(pwdata[13]),
    .B(\mem[8] [13]),
    .S(_1787_),
    .Z(_0816_));
 MUX2_X1 _4210_ (.A(pwdata[14]),
    .B(\mem[8] [14]),
    .S(_1787_),
    .Z(_0817_));
 MUX2_X1 _4211_ (.A(pwdata[15]),
    .B(\mem[8] [15]),
    .S(_1787_),
    .Z(_0818_));
 MUX2_X1 _4212_ (.A(pwdata[16]),
    .B(\mem[8] [16]),
    .S(_1787_),
    .Z(_0819_));
 MUX2_X1 _4213_ (.A(pwdata[17]),
    .B(\mem[8] [17]),
    .S(_1787_),
    .Z(_0820_));
 MUX2_X1 _4214_ (.A(pwdata[18]),
    .B(\mem[8] [18]),
    .S(_1787_),
    .Z(_0821_));
 MUX2_X1 _4215_ (.A(pwdata[19]),
    .B(\mem[8] [19]),
    .S(_1787_),
    .Z(_0822_));
 MUX2_X1 _4216_ (.A(pwdata[20]),
    .B(\mem[8] [20]),
    .S(_1787_),
    .Z(_0823_));
 MUX2_X1 _4217_ (.A(pwdata[21]),
    .B(\mem[8] [21]),
    .S(_1787_),
    .Z(_0824_));
 MUX2_X1 _4218_ (.A(pwdata[22]),
    .B(\mem[8] [22]),
    .S(_1787_),
    .Z(_0825_));
 MUX2_X1 _4219_ (.A(pwdata[23]),
    .B(\mem[8] [23]),
    .S(_1787_),
    .Z(_0826_));
 MUX2_X1 _4220_ (.A(pwdata[24]),
    .B(\mem[8] [24]),
    .S(_1787_),
    .Z(_0827_));
 MUX2_X1 _4221_ (.A(pwdata[25]),
    .B(\mem[8] [25]),
    .S(_1787_),
    .Z(_0828_));
 MUX2_X1 _4222_ (.A(pwdata[26]),
    .B(\mem[8] [26]),
    .S(_1787_),
    .Z(_0829_));
 MUX2_X1 _4223_ (.A(pwdata[27]),
    .B(\mem[8] [27]),
    .S(_1787_),
    .Z(_0830_));
 MUX2_X1 _4224_ (.A(pwdata[28]),
    .B(\mem[8] [28]),
    .S(_1787_),
    .Z(_0831_));
 MUX2_X1 _4225_ (.A(pwdata[29]),
    .B(\mem[8] [29]),
    .S(_1787_),
    .Z(_0832_));
 MUX2_X1 _4226_ (.A(pwdata[30]),
    .B(\mem[8] [30]),
    .S(_1787_),
    .Z(_0833_));
 MUX2_X1 _4227_ (.A(pwdata[31]),
    .B(\mem[8] [31]),
    .S(_1787_),
    .Z(_0834_));
 NAND2_X4 _4228_ (.A1(_1090_),
    .A2(_1138_),
    .ZN(_1788_));
 MUX2_X1 _4229_ (.A(pwdata[0]),
    .B(\mem[5] [0]),
    .S(_1788_),
    .Z(_0835_));
 MUX2_X1 _4230_ (.A(pwdata[1]),
    .B(\mem[5] [1]),
    .S(_1788_),
    .Z(_0836_));
 MUX2_X1 _4231_ (.A(pwdata[2]),
    .B(\mem[5] [2]),
    .S(_1788_),
    .Z(_0837_));
 MUX2_X1 _4232_ (.A(pwdata[3]),
    .B(\mem[5] [3]),
    .S(_1788_),
    .Z(_0838_));
 MUX2_X1 _4233_ (.A(pwdata[4]),
    .B(\mem[5] [4]),
    .S(_1788_),
    .Z(_0839_));
 MUX2_X1 _4234_ (.A(pwdata[5]),
    .B(\mem[5] [5]),
    .S(_1788_),
    .Z(_0840_));
 MUX2_X1 _4235_ (.A(pwdata[6]),
    .B(\mem[5] [6]),
    .S(_1788_),
    .Z(_0841_));
 MUX2_X1 _4236_ (.A(pwdata[7]),
    .B(\mem[5] [7]),
    .S(_1788_),
    .Z(_0842_));
 MUX2_X1 _4237_ (.A(pwdata[8]),
    .B(\mem[5] [8]),
    .S(_1788_),
    .Z(_0843_));
 MUX2_X1 _4238_ (.A(pwdata[9]),
    .B(\mem[5] [9]),
    .S(_1788_),
    .Z(_0844_));
 MUX2_X1 _4239_ (.A(pwdata[10]),
    .B(\mem[5] [10]),
    .S(_1788_),
    .Z(_0845_));
 MUX2_X1 _4240_ (.A(pwdata[11]),
    .B(\mem[5] [11]),
    .S(_1788_),
    .Z(_0846_));
 MUX2_X1 _4241_ (.A(pwdata[12]),
    .B(\mem[5] [12]),
    .S(_1788_),
    .Z(_0847_));
 MUX2_X1 _4242_ (.A(pwdata[13]),
    .B(\mem[5] [13]),
    .S(_1788_),
    .Z(_0848_));
 MUX2_X1 _4243_ (.A(pwdata[14]),
    .B(\mem[5] [14]),
    .S(_1788_),
    .Z(_0849_));
 MUX2_X1 _4244_ (.A(pwdata[15]),
    .B(\mem[5] [15]),
    .S(_1788_),
    .Z(_0850_));
 MUX2_X1 _4245_ (.A(pwdata[16]),
    .B(\mem[5] [16]),
    .S(_1788_),
    .Z(_0851_));
 MUX2_X1 _4246_ (.A(pwdata[17]),
    .B(\mem[5] [17]),
    .S(_1788_),
    .Z(_0852_));
 MUX2_X1 _4247_ (.A(pwdata[18]),
    .B(\mem[5] [18]),
    .S(_1788_),
    .Z(_0853_));
 MUX2_X1 _4248_ (.A(pwdata[19]),
    .B(\mem[5] [19]),
    .S(_1788_),
    .Z(_0854_));
 MUX2_X1 _4249_ (.A(pwdata[20]),
    .B(\mem[5] [20]),
    .S(_1788_),
    .Z(_0855_));
 MUX2_X1 _4250_ (.A(pwdata[21]),
    .B(\mem[5] [21]),
    .S(_1788_),
    .Z(_0856_));
 MUX2_X1 _4251_ (.A(pwdata[22]),
    .B(\mem[5] [22]),
    .S(_1788_),
    .Z(_0857_));
 MUX2_X1 _4252_ (.A(pwdata[23]),
    .B(\mem[5] [23]),
    .S(_1788_),
    .Z(_0858_));
 MUX2_X1 _4253_ (.A(pwdata[24]),
    .B(\mem[5] [24]),
    .S(_1788_),
    .Z(_0859_));
 MUX2_X1 _4254_ (.A(pwdata[25]),
    .B(\mem[5] [25]),
    .S(_1788_),
    .Z(_0860_));
 MUX2_X1 _4255_ (.A(pwdata[26]),
    .B(\mem[5] [26]),
    .S(_1788_),
    .Z(_0861_));
 MUX2_X1 _4256_ (.A(pwdata[27]),
    .B(\mem[5] [27]),
    .S(_1788_),
    .Z(_0862_));
 MUX2_X1 _4257_ (.A(pwdata[28]),
    .B(\mem[5] [28]),
    .S(_1788_),
    .Z(_0863_));
 MUX2_X1 _4258_ (.A(pwdata[29]),
    .B(\mem[5] [29]),
    .S(_1788_),
    .Z(_0864_));
 MUX2_X1 _4259_ (.A(pwdata[30]),
    .B(\mem[5] [30]),
    .S(_1788_),
    .Z(_0865_));
 MUX2_X1 _4260_ (.A(pwdata[31]),
    .B(\mem[5] [31]),
    .S(_1788_),
    .Z(_0866_));
 NAND2_X4 _4261_ (.A1(net2),
    .A2(net46),
    .ZN(_1789_));
 MUX2_X1 _4262_ (.A(pwdata[0]),
    .B(\mem[0] [0]),
    .S(_1789_),
    .Z(_0867_));
 MUX2_X1 _4263_ (.A(pwdata[1]),
    .B(\mem[0] [1]),
    .S(_1789_),
    .Z(_0868_));
 MUX2_X1 _4264_ (.A(pwdata[2]),
    .B(\mem[0] [2]),
    .S(_1789_),
    .Z(_0869_));
 MUX2_X1 _4265_ (.A(pwdata[3]),
    .B(\mem[0] [3]),
    .S(_1789_),
    .Z(_0870_));
 MUX2_X1 _4266_ (.A(pwdata[4]),
    .B(\mem[0] [4]),
    .S(_1789_),
    .Z(_0871_));
 MUX2_X1 _4267_ (.A(pwdata[5]),
    .B(\mem[0] [5]),
    .S(_1789_),
    .Z(_0872_));
 MUX2_X1 _4268_ (.A(pwdata[6]),
    .B(\mem[0] [6]),
    .S(_1789_),
    .Z(_0873_));
 MUX2_X1 _4269_ (.A(pwdata[7]),
    .B(\mem[0] [7]),
    .S(_1789_),
    .Z(_0874_));
 MUX2_X1 _4270_ (.A(pwdata[8]),
    .B(\mem[0] [8]),
    .S(_1789_),
    .Z(_0875_));
 MUX2_X1 _4271_ (.A(pwdata[9]),
    .B(\mem[0] [9]),
    .S(_1789_),
    .Z(_0876_));
 MUX2_X1 _4272_ (.A(pwdata[10]),
    .B(\mem[0] [10]),
    .S(_1789_),
    .Z(_0877_));
 MUX2_X1 _4273_ (.A(pwdata[11]),
    .B(\mem[0] [11]),
    .S(_1789_),
    .Z(_0878_));
 MUX2_X1 _4274_ (.A(pwdata[12]),
    .B(\mem[0] [12]),
    .S(_1789_),
    .Z(_0879_));
 MUX2_X1 _4275_ (.A(pwdata[13]),
    .B(\mem[0] [13]),
    .S(_1789_),
    .Z(_0880_));
 MUX2_X1 _4276_ (.A(pwdata[14]),
    .B(\mem[0] [14]),
    .S(_1789_),
    .Z(_0881_));
 MUX2_X1 _4277_ (.A(pwdata[15]),
    .B(\mem[0] [15]),
    .S(_1789_),
    .Z(_0882_));
 MUX2_X1 _4278_ (.A(pwdata[16]),
    .B(\mem[0] [16]),
    .S(_1789_),
    .Z(_0883_));
 MUX2_X1 _4279_ (.A(pwdata[17]),
    .B(\mem[0] [17]),
    .S(_1789_),
    .Z(_0884_));
 MUX2_X1 _4280_ (.A(pwdata[18]),
    .B(\mem[0] [18]),
    .S(_1789_),
    .Z(_0885_));
 MUX2_X1 _4281_ (.A(pwdata[19]),
    .B(\mem[0] [19]),
    .S(_1789_),
    .Z(_0886_));
 MUX2_X1 _4282_ (.A(pwdata[20]),
    .B(\mem[0] [20]),
    .S(_1789_),
    .Z(_0887_));
 MUX2_X1 _4283_ (.A(pwdata[21]),
    .B(\mem[0] [21]),
    .S(_1789_),
    .Z(_0888_));
 MUX2_X1 _4284_ (.A(pwdata[22]),
    .B(\mem[0] [22]),
    .S(_1789_),
    .Z(_0889_));
 MUX2_X1 _4285_ (.A(pwdata[23]),
    .B(\mem[0] [23]),
    .S(_1789_),
    .Z(_0890_));
 MUX2_X1 _4286_ (.A(pwdata[24]),
    .B(\mem[0] [24]),
    .S(_1789_),
    .Z(_0891_));
 MUX2_X1 _4287_ (.A(pwdata[25]),
    .B(\mem[0] [25]),
    .S(_1789_),
    .Z(_0892_));
 MUX2_X1 _4288_ (.A(pwdata[26]),
    .B(\mem[0] [26]),
    .S(_1789_),
    .Z(_0893_));
 MUX2_X1 _4289_ (.A(pwdata[27]),
    .B(\mem[0] [27]),
    .S(_1789_),
    .Z(_0894_));
 MUX2_X1 _4290_ (.A(pwdata[28]),
    .B(\mem[0] [28]),
    .S(_1789_),
    .Z(_0895_));
 MUX2_X1 _4291_ (.A(pwdata[29]),
    .B(\mem[0] [29]),
    .S(_1789_),
    .Z(_0896_));
 MUX2_X1 _4292_ (.A(pwdata[30]),
    .B(\mem[0] [30]),
    .S(_1789_),
    .Z(_0897_));
 MUX2_X1 _4293_ (.A(pwdata[31]),
    .B(\mem[0] [31]),
    .S(_1789_),
    .Z(_0898_));
 NAND2_X4 _4294_ (.A1(net2),
    .A2(net41),
    .ZN(_1790_));
 MUX2_X1 _4295_ (.A(pwdata[0]),
    .B(\mem[4] [0]),
    .S(_1790_),
    .Z(_0899_));
 MUX2_X1 _4296_ (.A(pwdata[1]),
    .B(\mem[4] [1]),
    .S(_1790_),
    .Z(_0900_));
 MUX2_X1 _4297_ (.A(pwdata[2]),
    .B(\mem[4] [2]),
    .S(_1790_),
    .Z(_0901_));
 MUX2_X1 _4298_ (.A(pwdata[3]),
    .B(\mem[4] [3]),
    .S(_1790_),
    .Z(_0902_));
 MUX2_X1 _4299_ (.A(pwdata[4]),
    .B(\mem[4] [4]),
    .S(_1790_),
    .Z(_0903_));
 MUX2_X1 _4300_ (.A(pwdata[5]),
    .B(\mem[4] [5]),
    .S(_1790_),
    .Z(_0904_));
 MUX2_X1 _4301_ (.A(pwdata[6]),
    .B(\mem[4] [6]),
    .S(_1790_),
    .Z(_0905_));
 MUX2_X1 _4302_ (.A(pwdata[7]),
    .B(\mem[4] [7]),
    .S(_1790_),
    .Z(_0906_));
 MUX2_X1 _4303_ (.A(pwdata[8]),
    .B(\mem[4] [8]),
    .S(_1790_),
    .Z(_0907_));
 MUX2_X1 _4304_ (.A(pwdata[9]),
    .B(\mem[4] [9]),
    .S(_1790_),
    .Z(_0908_));
 MUX2_X1 _4305_ (.A(pwdata[10]),
    .B(\mem[4] [10]),
    .S(_1790_),
    .Z(_0909_));
 MUX2_X1 _4306_ (.A(pwdata[11]),
    .B(\mem[4] [11]),
    .S(_1790_),
    .Z(_0910_));
 MUX2_X1 _4307_ (.A(pwdata[12]),
    .B(\mem[4] [12]),
    .S(_1790_),
    .Z(_0911_));
 MUX2_X1 _4308_ (.A(pwdata[13]),
    .B(\mem[4] [13]),
    .S(_1790_),
    .Z(_0912_));
 MUX2_X1 _4309_ (.A(pwdata[14]),
    .B(\mem[4] [14]),
    .S(_1790_),
    .Z(_0913_));
 MUX2_X1 _4310_ (.A(pwdata[15]),
    .B(\mem[4] [15]),
    .S(_1790_),
    .Z(_0914_));
 MUX2_X1 _4311_ (.A(pwdata[16]),
    .B(\mem[4] [16]),
    .S(_1790_),
    .Z(_0915_));
 MUX2_X1 _4312_ (.A(pwdata[17]),
    .B(\mem[4] [17]),
    .S(_1790_),
    .Z(_0916_));
 MUX2_X1 _4313_ (.A(pwdata[18]),
    .B(\mem[4] [18]),
    .S(_1790_),
    .Z(_0917_));
 MUX2_X1 _4314_ (.A(pwdata[19]),
    .B(\mem[4] [19]),
    .S(_1790_),
    .Z(_0918_));
 MUX2_X1 _4315_ (.A(pwdata[20]),
    .B(\mem[4] [20]),
    .S(_1790_),
    .Z(_0919_));
 MUX2_X1 _4316_ (.A(pwdata[21]),
    .B(\mem[4] [21]),
    .S(_1790_),
    .Z(_0920_));
 MUX2_X1 _4317_ (.A(pwdata[22]),
    .B(\mem[4] [22]),
    .S(_1790_),
    .Z(_0921_));
 MUX2_X1 _4318_ (.A(pwdata[23]),
    .B(\mem[4] [23]),
    .S(_1790_),
    .Z(_0922_));
 MUX2_X1 _4319_ (.A(pwdata[24]),
    .B(\mem[4] [24]),
    .S(_1790_),
    .Z(_0923_));
 MUX2_X1 _4320_ (.A(pwdata[25]),
    .B(\mem[4] [25]),
    .S(_1790_),
    .Z(_0924_));
 MUX2_X1 _4321_ (.A(pwdata[26]),
    .B(\mem[4] [26]),
    .S(_1790_),
    .Z(_0925_));
 MUX2_X1 _4322_ (.A(pwdata[27]),
    .B(\mem[4] [27]),
    .S(_1790_),
    .Z(_0926_));
 MUX2_X1 _4323_ (.A(pwdata[28]),
    .B(\mem[4] [28]),
    .S(_1790_),
    .Z(_0927_));
 MUX2_X1 _4324_ (.A(pwdata[29]),
    .B(\mem[4] [29]),
    .S(_1790_),
    .Z(_0928_));
 MUX2_X1 _4325_ (.A(pwdata[30]),
    .B(\mem[4] [30]),
    .S(_1790_),
    .Z(_0929_));
 MUX2_X1 _4326_ (.A(pwdata[31]),
    .B(\mem[4] [31]),
    .S(_1790_),
    .Z(_0930_));
 NAND2_X4 _4327_ (.A1(net2),
    .A2(_1147_),
    .ZN(_1791_));
 MUX2_X1 _4328_ (.A(pwdata[0]),
    .B(\mem[6] [0]),
    .S(_1791_),
    .Z(_0931_));
 MUX2_X1 _4329_ (.A(pwdata[1]),
    .B(\mem[6] [1]),
    .S(_1791_),
    .Z(_0932_));
 MUX2_X1 _4330_ (.A(pwdata[2]),
    .B(\mem[6] [2]),
    .S(_1791_),
    .Z(_0933_));
 MUX2_X1 _4331_ (.A(pwdata[3]),
    .B(\mem[6] [3]),
    .S(_1791_),
    .Z(_0934_));
 MUX2_X1 _4332_ (.A(pwdata[4]),
    .B(\mem[6] [4]),
    .S(_1791_),
    .Z(_0935_));
 MUX2_X1 _4333_ (.A(pwdata[5]),
    .B(\mem[6] [5]),
    .S(_1791_),
    .Z(_0936_));
 MUX2_X1 _4334_ (.A(pwdata[6]),
    .B(\mem[6] [6]),
    .S(_1791_),
    .Z(_0937_));
 MUX2_X1 _4335_ (.A(pwdata[7]),
    .B(\mem[6] [7]),
    .S(_1791_),
    .Z(_0938_));
 MUX2_X1 _4336_ (.A(pwdata[8]),
    .B(\mem[6] [8]),
    .S(_1791_),
    .Z(_0939_));
 MUX2_X1 _4337_ (.A(pwdata[9]),
    .B(\mem[6] [9]),
    .S(_1791_),
    .Z(_0940_));
 MUX2_X1 _4338_ (.A(pwdata[10]),
    .B(\mem[6] [10]),
    .S(_1791_),
    .Z(_0941_));
 MUX2_X1 _4339_ (.A(pwdata[11]),
    .B(\mem[6] [11]),
    .S(_1791_),
    .Z(_0942_));
 MUX2_X1 _4340_ (.A(pwdata[12]),
    .B(\mem[6] [12]),
    .S(_1791_),
    .Z(_0943_));
 MUX2_X1 _4341_ (.A(pwdata[13]),
    .B(\mem[6] [13]),
    .S(_1791_),
    .Z(_0944_));
 MUX2_X1 _4342_ (.A(pwdata[14]),
    .B(\mem[6] [14]),
    .S(_1791_),
    .Z(_0945_));
 MUX2_X1 _4343_ (.A(pwdata[15]),
    .B(\mem[6] [15]),
    .S(_1791_),
    .Z(_0946_));
 MUX2_X1 _4344_ (.A(pwdata[16]),
    .B(\mem[6] [16]),
    .S(_1791_),
    .Z(_0947_));
 MUX2_X1 _4345_ (.A(pwdata[17]),
    .B(\mem[6] [17]),
    .S(_1791_),
    .Z(_0948_));
 MUX2_X1 _4346_ (.A(pwdata[18]),
    .B(\mem[6] [18]),
    .S(_1791_),
    .Z(_0949_));
 MUX2_X1 _4347_ (.A(pwdata[19]),
    .B(\mem[6] [19]),
    .S(_1791_),
    .Z(_0950_));
 MUX2_X1 _4348_ (.A(pwdata[20]),
    .B(\mem[6] [20]),
    .S(_1791_),
    .Z(_0951_));
 MUX2_X1 _4349_ (.A(pwdata[21]),
    .B(\mem[6] [21]),
    .S(_1791_),
    .Z(_0952_));
 MUX2_X1 _4350_ (.A(pwdata[22]),
    .B(\mem[6] [22]),
    .S(_1791_),
    .Z(_0953_));
 MUX2_X1 _4351_ (.A(pwdata[23]),
    .B(\mem[6] [23]),
    .S(_1791_),
    .Z(_0954_));
 MUX2_X1 _4352_ (.A(pwdata[24]),
    .B(\mem[6] [24]),
    .S(_1791_),
    .Z(_0955_));
 MUX2_X1 _4353_ (.A(pwdata[25]),
    .B(\mem[6] [25]),
    .S(_1791_),
    .Z(_0956_));
 MUX2_X1 _4354_ (.A(pwdata[26]),
    .B(\mem[6] [26]),
    .S(_1791_),
    .Z(_0957_));
 MUX2_X1 _4355_ (.A(pwdata[27]),
    .B(\mem[6] [27]),
    .S(_1791_),
    .Z(_0958_));
 MUX2_X1 _4356_ (.A(pwdata[28]),
    .B(\mem[6] [28]),
    .S(_1791_),
    .Z(_0959_));
 MUX2_X1 _4357_ (.A(pwdata[29]),
    .B(\mem[6] [29]),
    .S(_1791_),
    .Z(_0960_));
 MUX2_X1 _4358_ (.A(pwdata[30]),
    .B(\mem[6] [30]),
    .S(_1791_),
    .Z(_0961_));
 MUX2_X1 _4359_ (.A(pwdata[31]),
    .B(\mem[6] [31]),
    .S(_1791_),
    .Z(_0962_));
 NAND2_X4 _4360_ (.A1(net2),
    .A2(net31),
    .ZN(_1792_));
 MUX2_X1 _4361_ (.A(pwdata[0]),
    .B(\mem[13] [0]),
    .S(_1792_),
    .Z(_0963_));
 MUX2_X1 _4362_ (.A(pwdata[1]),
    .B(\mem[13] [1]),
    .S(_1792_),
    .Z(_0964_));
 MUX2_X1 _4363_ (.A(pwdata[2]),
    .B(\mem[13] [2]),
    .S(_1792_),
    .Z(_0965_));
 MUX2_X1 _4364_ (.A(pwdata[3]),
    .B(\mem[13] [3]),
    .S(_1792_),
    .Z(_0966_));
 MUX2_X1 _4365_ (.A(pwdata[4]),
    .B(\mem[13] [4]),
    .S(_1792_),
    .Z(_0967_));
 MUX2_X1 _4366_ (.A(pwdata[5]),
    .B(\mem[13] [5]),
    .S(_1792_),
    .Z(_0968_));
 MUX2_X1 _4367_ (.A(pwdata[6]),
    .B(\mem[13] [6]),
    .S(_1792_),
    .Z(_0969_));
 MUX2_X1 _4368_ (.A(pwdata[7]),
    .B(\mem[13] [7]),
    .S(_1792_),
    .Z(_0970_));
 MUX2_X1 _4369_ (.A(pwdata[8]),
    .B(\mem[13] [8]),
    .S(_1792_),
    .Z(_0971_));
 MUX2_X1 _4370_ (.A(pwdata[9]),
    .B(\mem[13] [9]),
    .S(_1792_),
    .Z(_0972_));
 MUX2_X1 _4371_ (.A(pwdata[10]),
    .B(\mem[13] [10]),
    .S(_1792_),
    .Z(_0973_));
 MUX2_X1 _4372_ (.A(pwdata[11]),
    .B(\mem[13] [11]),
    .S(_1792_),
    .Z(_0974_));
 MUX2_X1 _4373_ (.A(pwdata[12]),
    .B(\mem[13] [12]),
    .S(_1792_),
    .Z(_0975_));
 MUX2_X1 _4374_ (.A(pwdata[13]),
    .B(\mem[13] [13]),
    .S(_1792_),
    .Z(_0976_));
 MUX2_X1 _4375_ (.A(pwdata[14]),
    .B(\mem[13] [14]),
    .S(_1792_),
    .Z(_0977_));
 MUX2_X1 _4376_ (.A(pwdata[15]),
    .B(\mem[13] [15]),
    .S(_1792_),
    .Z(_0978_));
 MUX2_X1 _4377_ (.A(pwdata[16]),
    .B(\mem[13] [16]),
    .S(_1792_),
    .Z(_0979_));
 MUX2_X1 _4378_ (.A(pwdata[17]),
    .B(\mem[13] [17]),
    .S(_1792_),
    .Z(_0980_));
 MUX2_X1 _4379_ (.A(pwdata[18]),
    .B(\mem[13] [18]),
    .S(_1792_),
    .Z(_0981_));
 MUX2_X1 _4380_ (.A(pwdata[19]),
    .B(\mem[13] [19]),
    .S(_1792_),
    .Z(_0982_));
 MUX2_X1 _4381_ (.A(pwdata[20]),
    .B(\mem[13] [20]),
    .S(_1792_),
    .Z(_0983_));
 MUX2_X1 _4382_ (.A(pwdata[21]),
    .B(\mem[13] [21]),
    .S(_1792_),
    .Z(_0984_));
 MUX2_X1 _4383_ (.A(pwdata[22]),
    .B(\mem[13] [22]),
    .S(_1792_),
    .Z(_0985_));
 MUX2_X1 _4384_ (.A(pwdata[23]),
    .B(\mem[13] [23]),
    .S(_1792_),
    .Z(_0986_));
 MUX2_X1 _4385_ (.A(pwdata[24]),
    .B(\mem[13] [24]),
    .S(_1792_),
    .Z(_0987_));
 MUX2_X1 _4386_ (.A(pwdata[25]),
    .B(\mem[13] [25]),
    .S(_1792_),
    .Z(_0988_));
 MUX2_X1 _4387_ (.A(pwdata[26]),
    .B(\mem[13] [26]),
    .S(_1792_),
    .Z(_0989_));
 MUX2_X1 _4388_ (.A(pwdata[27]),
    .B(\mem[13] [27]),
    .S(_1792_),
    .Z(_0990_));
 MUX2_X1 _4389_ (.A(pwdata[28]),
    .B(\mem[13] [28]),
    .S(_1792_),
    .Z(_0991_));
 MUX2_X1 _4390_ (.A(pwdata[29]),
    .B(\mem[13] [29]),
    .S(_1792_),
    .Z(_0992_));
 MUX2_X1 _4391_ (.A(pwdata[30]),
    .B(\mem[13] [30]),
    .S(_1792_),
    .Z(_0993_));
 MUX2_X1 _4392_ (.A(pwdata[31]),
    .B(\mem[13] [31]),
    .S(_1792_),
    .Z(_0994_));
 NAND2_X4 _4393_ (.A1(net2),
    .A2(net29),
    .ZN(_1793_));
 MUX2_X1 _4394_ (.A(pwdata[0]),
    .B(\mem[14] [0]),
    .S(_1793_),
    .Z(_0995_));
 MUX2_X1 _4395_ (.A(pwdata[1]),
    .B(\mem[14] [1]),
    .S(_1793_),
    .Z(_0996_));
 MUX2_X1 _4396_ (.A(pwdata[2]),
    .B(\mem[14] [2]),
    .S(_1793_),
    .Z(_0997_));
 MUX2_X1 _4397_ (.A(pwdata[3]),
    .B(\mem[14] [3]),
    .S(_1793_),
    .Z(_0998_));
 MUX2_X1 _4398_ (.A(pwdata[4]),
    .B(\mem[14] [4]),
    .S(_1793_),
    .Z(_0999_));
 MUX2_X1 _4399_ (.A(pwdata[5]),
    .B(\mem[14] [5]),
    .S(_1793_),
    .Z(_1000_));
 MUX2_X1 _4400_ (.A(pwdata[6]),
    .B(\mem[14] [6]),
    .S(_1793_),
    .Z(_1001_));
 MUX2_X1 _4401_ (.A(pwdata[7]),
    .B(\mem[14] [7]),
    .S(_1793_),
    .Z(_1002_));
 MUX2_X1 _4402_ (.A(pwdata[8]),
    .B(\mem[14] [8]),
    .S(_1793_),
    .Z(_1003_));
 MUX2_X1 _4403_ (.A(pwdata[9]),
    .B(\mem[14] [9]),
    .S(_1793_),
    .Z(_1004_));
 MUX2_X1 _4404_ (.A(pwdata[10]),
    .B(\mem[14] [10]),
    .S(_1793_),
    .Z(_1005_));
 MUX2_X1 _4405_ (.A(pwdata[11]),
    .B(\mem[14] [11]),
    .S(_1793_),
    .Z(_1006_));
 MUX2_X1 _4406_ (.A(pwdata[12]),
    .B(\mem[14] [12]),
    .S(_1793_),
    .Z(_1007_));
 MUX2_X1 _4407_ (.A(pwdata[13]),
    .B(\mem[14] [13]),
    .S(_1793_),
    .Z(_1008_));
 MUX2_X1 _4408_ (.A(pwdata[14]),
    .B(\mem[14] [14]),
    .S(_1793_),
    .Z(_1009_));
 MUX2_X1 _4409_ (.A(pwdata[15]),
    .B(\mem[14] [15]),
    .S(_1793_),
    .Z(_1010_));
 MUX2_X1 _4410_ (.A(pwdata[16]),
    .B(\mem[14] [16]),
    .S(_1793_),
    .Z(_1011_));
 MUX2_X1 _4411_ (.A(pwdata[17]),
    .B(\mem[14] [17]),
    .S(_1793_),
    .Z(_1012_));
 MUX2_X1 _4412_ (.A(pwdata[18]),
    .B(\mem[14] [18]),
    .S(_1793_),
    .Z(_1013_));
 MUX2_X1 _4413_ (.A(pwdata[19]),
    .B(\mem[14] [19]),
    .S(_1793_),
    .Z(_1014_));
 MUX2_X1 _4414_ (.A(pwdata[20]),
    .B(\mem[14] [20]),
    .S(_1793_),
    .Z(_1015_));
 MUX2_X1 _4415_ (.A(pwdata[21]),
    .B(\mem[14] [21]),
    .S(_1793_),
    .Z(_1016_));
 MUX2_X1 _4416_ (.A(pwdata[22]),
    .B(\mem[14] [22]),
    .S(_1793_),
    .Z(_1017_));
 MUX2_X1 _4417_ (.A(pwdata[23]),
    .B(\mem[14] [23]),
    .S(_1793_),
    .Z(_1018_));
 MUX2_X1 _4418_ (.A(pwdata[24]),
    .B(\mem[14] [24]),
    .S(_1793_),
    .Z(_1019_));
 MUX2_X1 _4419_ (.A(pwdata[25]),
    .B(\mem[14] [25]),
    .S(_1793_),
    .Z(_1020_));
 MUX2_X1 _4420_ (.A(pwdata[26]),
    .B(\mem[14] [26]),
    .S(_1793_),
    .Z(_1021_));
 MUX2_X1 _4421_ (.A(pwdata[27]),
    .B(\mem[14] [27]),
    .S(_1793_),
    .Z(_1022_));
 MUX2_X1 _4422_ (.A(pwdata[28]),
    .B(\mem[14] [28]),
    .S(_1793_),
    .Z(_1023_));
 MUX2_X1 _4423_ (.A(pwdata[29]),
    .B(\mem[14] [29]),
    .S(_1793_),
    .Z(_1024_));
 MUX2_X1 _4424_ (.A(pwdata[30]),
    .B(\mem[14] [30]),
    .S(_1793_),
    .Z(_1025_));
 MUX2_X1 _4425_ (.A(pwdata[31]),
    .B(\mem[14] [31]),
    .S(_1793_),
    .Z(_1026_));
 NAND2_X4 _4426_ (.A1(net2),
    .A2(net38),
    .ZN(_1794_));
 MUX2_X1 _4427_ (.A(pwdata[0]),
    .B(\mem[11] [0]),
    .S(_1794_),
    .Z(_1027_));
 MUX2_X1 _4428_ (.A(pwdata[1]),
    .B(\mem[11] [1]),
    .S(_1794_),
    .Z(_1028_));
 MUX2_X1 _4429_ (.A(pwdata[2]),
    .B(\mem[11] [2]),
    .S(_1794_),
    .Z(_1029_));
 MUX2_X1 _4430_ (.A(pwdata[3]),
    .B(\mem[11] [3]),
    .S(_1794_),
    .Z(_1030_));
 MUX2_X1 _4431_ (.A(pwdata[4]),
    .B(\mem[11] [4]),
    .S(_1794_),
    .Z(_1031_));
 MUX2_X1 _4432_ (.A(pwdata[5]),
    .B(\mem[11] [5]),
    .S(_1794_),
    .Z(_1032_));
 MUX2_X1 _4433_ (.A(pwdata[6]),
    .B(\mem[11] [6]),
    .S(_1794_),
    .Z(_1033_));
 MUX2_X1 _4434_ (.A(pwdata[7]),
    .B(\mem[11] [7]),
    .S(_1794_),
    .Z(_1034_));
 MUX2_X1 _4435_ (.A(pwdata[8]),
    .B(\mem[11] [8]),
    .S(_1794_),
    .Z(_1035_));
 MUX2_X1 _4436_ (.A(pwdata[9]),
    .B(\mem[11] [9]),
    .S(_1794_),
    .Z(_1036_));
 MUX2_X1 _4437_ (.A(pwdata[10]),
    .B(\mem[11] [10]),
    .S(_1794_),
    .Z(_1037_));
 MUX2_X1 _4438_ (.A(pwdata[11]),
    .B(\mem[11] [11]),
    .S(_1794_),
    .Z(_1038_));
 MUX2_X1 _4439_ (.A(pwdata[12]),
    .B(\mem[11] [12]),
    .S(_1794_),
    .Z(_1039_));
 MUX2_X1 _4440_ (.A(pwdata[13]),
    .B(\mem[11] [13]),
    .S(_1794_),
    .Z(_1040_));
 MUX2_X1 _4441_ (.A(pwdata[14]),
    .B(\mem[11] [14]),
    .S(_1794_),
    .Z(_1041_));
 MUX2_X1 _4442_ (.A(pwdata[15]),
    .B(\mem[11] [15]),
    .S(_1794_),
    .Z(_1042_));
 MUX2_X1 _4443_ (.A(pwdata[16]),
    .B(\mem[11] [16]),
    .S(_1794_),
    .Z(_1043_));
 MUX2_X1 _4444_ (.A(pwdata[17]),
    .B(\mem[11] [17]),
    .S(_1794_),
    .Z(_1044_));
 MUX2_X1 _4445_ (.A(pwdata[18]),
    .B(\mem[11] [18]),
    .S(_1794_),
    .Z(_1045_));
 MUX2_X1 _4446_ (.A(pwdata[19]),
    .B(\mem[11] [19]),
    .S(_1794_),
    .Z(_1046_));
 MUX2_X1 _4447_ (.A(pwdata[20]),
    .B(\mem[11] [20]),
    .S(_1794_),
    .Z(_1047_));
 MUX2_X1 _4448_ (.A(pwdata[21]),
    .B(\mem[11] [21]),
    .S(_1794_),
    .Z(_1048_));
 MUX2_X1 _4449_ (.A(pwdata[22]),
    .B(\mem[11] [22]),
    .S(_1794_),
    .Z(_1049_));
 MUX2_X1 _4450_ (.A(pwdata[23]),
    .B(\mem[11] [23]),
    .S(_1794_),
    .Z(_1050_));
 MUX2_X1 _4451_ (.A(pwdata[24]),
    .B(\mem[11] [24]),
    .S(_1794_),
    .Z(_1051_));
 MUX2_X1 _4452_ (.A(pwdata[25]),
    .B(\mem[11] [25]),
    .S(_1794_),
    .Z(_1052_));
 MUX2_X1 _4453_ (.A(pwdata[26]),
    .B(\mem[11] [26]),
    .S(_1794_),
    .Z(_1053_));
 MUX2_X1 _4454_ (.A(pwdata[27]),
    .B(\mem[11] [27]),
    .S(_1794_),
    .Z(_1054_));
 MUX2_X1 _4455_ (.A(pwdata[28]),
    .B(\mem[11] [28]),
    .S(_1794_),
    .Z(_1055_));
 MUX2_X1 _4456_ (.A(pwdata[29]),
    .B(\mem[11] [29]),
    .S(_1794_),
    .Z(_1056_));
 MUX2_X1 _4457_ (.A(pwdata[30]),
    .B(\mem[11] [30]),
    .S(_1794_),
    .Z(_1057_));
 MUX2_X1 _4458_ (.A(pwdata[31]),
    .B(\mem[11] [31]),
    .S(_1794_),
    .Z(_1058_));
 OAI22_X1 _4459_ (.A1(present_state[1]),
    .A2(present_state[0]),
    .B1(penable),
    .B2(_1082_),
    .ZN(next_state[0]));
 NOR2_X1 _4460_ (.A1(present_state[1]),
    .A2(_0001_),
    .ZN(_1795_));
 AOI22_X1 _4461_ (.A1(penable),
    .A2(_2855_[0]),
    .B1(_1795_),
    .B2(pselx),
    .ZN(_1796_));
 INV_X1 _4462_ (.A(_1796_),
    .ZN(next_state[1]));
 INV_X1 _4463_ (.A(prdata[1]),
    .ZN(_1059_));
 INV_X1 _4464_ (.A(prdata[2]),
    .ZN(_1060_));
 INV_X1 _4465_ (.A(prdata[4]),
    .ZN(_1061_));
 INV_X1 _4466_ (.A(prdata[12]),
    .ZN(_1062_));
 INV_X1 _4467_ (.A(prdata[19]),
    .ZN(_1063_));
 INV_X1 _4468_ (.A(prdata[20]),
    .ZN(_1064_));
 INV_X1 _4469_ (.A(prdata[25]),
    .ZN(_1065_));
 INV_X1 _4470_ (.A(prdata[26]),
    .ZN(_1066_));
 INV_X1 _4471_ (.A(prdata[27]),
    .ZN(_1067_));
 INV_X1 _4472_ (.A(pslverr),
    .ZN(_1068_));
 INV_X2 _4473_ (.A(paddr[4]),
    .ZN(_1069_));
 INV_X2 _4474_ (.A(paddr[3]),
    .ZN(_1070_));
 INV_X2 _4475_ (.A(paddr[2]),
    .ZN(_1071_));
 INV_X2 _4476_ (.A(paddr[1]),
    .ZN(_1072_));
 INV_X2 _4477_ (.A(paddr[0]),
    .ZN(_1073_));
 INV_X1 _4478_ (.A(pwrite),
    .ZN(_1074_));
 NAND2_X4 _4479_ (.A1(paddr[3]),
    .A2(paddr[2]),
    .ZN(_1075_));
 OR2_X2 _4480_ (.A1(paddr[1]),
    .A2(paddr[0]),
    .ZN(_1076_));
 NOR3_X4 _4481_ (.A1(paddr[4]),
    .A2(_1075_),
    .A3(_1076_),
    .ZN(_1077_));
 NOR3_X1 _4482_ (.A1(paddr[5]),
    .A2(paddr[6]),
    .A3(paddr[7]),
    .ZN(_1078_));
 NOR4_X1 _4483_ (.A1(paddr[12]),
    .A2(paddr[13]),
    .A3(paddr[14]),
    .A4(paddr[15]),
    .ZN(_1079_));
 NOR4_X1 _4484_ (.A1(paddr[8]),
    .A2(paddr[9]),
    .A3(paddr[10]),
    .A4(paddr[11]),
    .ZN(_1080_));
 NAND3_X2 _4485_ (.A1(_1078_),
    .A2(_1079_),
    .A3(_1080_),
    .ZN(_1081_));
 NOR2_X2 _4486_ (.A1(present_state[0]),
    .A2(net71),
    .ZN(_2855_[0]));
 INV_X1 _4487_ (.A(_2855_[0]),
    .ZN(_1082_));
 NAND3_X1 _4488_ (.A1(pwrite),
    .A2(penable),
    .A3(_2855_[0]),
    .ZN(_1083_));
 NOR4_X2 _4489_ (.A1(paddr[20]),
    .A2(paddr[21]),
    .A3(paddr[22]),
    .A4(paddr[23]),
    .ZN(_1084_));
 NOR4_X1 _4490_ (.A1(paddr[16]),
    .A2(paddr[17]),
    .A3(paddr[18]),
    .A4(paddr[19]),
    .ZN(_1085_));
 NOR4_X1 _4491_ (.A1(paddr[28]),
    .A2(paddr[29]),
    .A3(paddr[30]),
    .A4(paddr[31]),
    .ZN(_1086_));
 NOR4_X1 _4492_ (.A1(paddr[24]),
    .A2(paddr[25]),
    .A3(paddr[26]),
    .A4(paddr[27]),
    .ZN(_1087_));
 NAND4_X1 _4493_ (.A1(_1084_),
    .A2(_1085_),
    .A3(_1086_),
    .A4(_1087_),
    .ZN(_1088_));
 NOR3_X1 _4494_ (.A1(_1081_),
    .A2(_1083_),
    .A3(_1088_),
    .ZN(_1089_));
 AND2_X4 _4495_ (.A1(prst_n),
    .A2(_1089_),
    .ZN(_1090_));
 NAND2_X4 _4496_ (.A1(net14),
    .A2(net2),
    .ZN(_1091_));
 MUX2_X1 _4497_ (.A(pwdata[0]),
    .B(\mem[12] [0]),
    .S(_1091_),
    .Z(_0002_));
 MUX2_X1 _4498_ (.A(pwdata[1]),
    .B(\mem[12] [1]),
    .S(_1091_),
    .Z(_0003_));
 MUX2_X1 _4499_ (.A(pwdata[2]),
    .B(\mem[12] [2]),
    .S(net1),
    .Z(_0004_));
 MUX2_X1 _4500_ (.A(pwdata[3]),
    .B(\mem[12] [3]),
    .S(net1),
    .Z(_0005_));
 MUX2_X1 _4501_ (.A(pwdata[4]),
    .B(\mem[12] [4]),
    .S(_1091_),
    .Z(_0006_));
 MUX2_X1 _4502_ (.A(pwdata[5]),
    .B(\mem[12] [5]),
    .S(net1),
    .Z(_0007_));
 MUX2_X1 _4503_ (.A(pwdata[6]),
    .B(\mem[12] [6]),
    .S(net1),
    .Z(_0008_));
 MUX2_X1 _4504_ (.A(pwdata[7]),
    .B(\mem[12] [7]),
    .S(_1091_),
    .Z(_0009_));
 MUX2_X1 _4505_ (.A(pwdata[8]),
    .B(\mem[12] [8]),
    .S(_1091_),
    .Z(_0010_));
 MUX2_X1 _4506_ (.A(pwdata[9]),
    .B(\mem[12] [9]),
    .S(net1),
    .Z(_0011_));
 MUX2_X1 _4507_ (.A(pwdata[10]),
    .B(\mem[12] [10]),
    .S(_1091_),
    .Z(_0012_));
 MUX2_X1 _4508_ (.A(pwdata[11]),
    .B(\mem[12] [11]),
    .S(net1),
    .Z(_0013_));
 MUX2_X1 _4509_ (.A(pwdata[12]),
    .B(\mem[12] [12]),
    .S(net1),
    .Z(_0014_));
 MUX2_X1 _4510_ (.A(pwdata[13]),
    .B(\mem[12] [13]),
    .S(_1091_),
    .Z(_0015_));
 MUX2_X1 _4511_ (.A(pwdata[14]),
    .B(\mem[12] [14]),
    .S(_1091_),
    .Z(_0016_));
 MUX2_X1 _4512_ (.A(pwdata[15]),
    .B(\mem[12] [15]),
    .S(_1091_),
    .Z(_0017_));
 MUX2_X1 _4513_ (.A(pwdata[16]),
    .B(\mem[12] [16]),
    .S(net1),
    .Z(_0018_));
 MUX2_X1 _4514_ (.A(pwdata[17]),
    .B(\mem[12] [17]),
    .S(net1),
    .Z(_0019_));
 MUX2_X1 _4515_ (.A(pwdata[18]),
    .B(\mem[12] [18]),
    .S(net1),
    .Z(_0020_));
 MUX2_X1 _4516_ (.A(pwdata[19]),
    .B(\mem[12] [19]),
    .S(net1),
    .Z(_0021_));
 MUX2_X1 _4517_ (.A(pwdata[20]),
    .B(\mem[12] [20]),
    .S(_1091_),
    .Z(_0022_));
 MUX2_X1 _4518_ (.A(pwdata[21]),
    .B(\mem[12] [21]),
    .S(net1),
    .Z(_0023_));
 MUX2_X1 _4519_ (.A(pwdata[22]),
    .B(\mem[12] [22]),
    .S(net1),
    .Z(_0024_));
 MUX2_X1 _4520_ (.A(pwdata[23]),
    .B(\mem[12] [23]),
    .S(net1),
    .Z(_0025_));
 MUX2_X1 _4521_ (.A(pwdata[24]),
    .B(\mem[12] [24]),
    .S(net1),
    .Z(_0026_));
 MUX2_X1 _4522_ (.A(pwdata[25]),
    .B(\mem[12] [25]),
    .S(_1091_),
    .Z(_0027_));
 MUX2_X1 _4523_ (.A(pwdata[26]),
    .B(\mem[12] [26]),
    .S(net1),
    .Z(_0028_));
 MUX2_X1 _4524_ (.A(pwdata[27]),
    .B(\mem[12] [27]),
    .S(net1),
    .Z(_0029_));
 MUX2_X1 _4525_ (.A(pwdata[28]),
    .B(\mem[12] [28]),
    .S(_1091_),
    .Z(_0030_));
 MUX2_X1 _4526_ (.A(pwdata[29]),
    .B(\mem[12] [29]),
    .S(_1091_),
    .Z(_0031_));
 MUX2_X1 _4527_ (.A(pwdata[30]),
    .B(\mem[12] [30]),
    .S(_1091_),
    .Z(_0032_));
 MUX2_X1 _4528_ (.A(pwdata[31]),
    .B(\mem[12] [31]),
    .S(_1091_),
    .Z(_0033_));
 NAND2_X4 _4529_ (.A1(paddr[1]),
    .A2(paddr[0]),
    .ZN(_1092_));
 NOR3_X4 _4530_ (.A1(paddr[4]),
    .A2(_1075_),
    .A3(_1092_),
    .ZN(_1093_));
 NAND2_X4 _4531_ (.A1(_1090_),
    .A2(_1093_),
    .ZN(_1094_));
 MUX2_X1 _4532_ (.A(pwdata[0]),
    .B(\mem[15] [0]),
    .S(_1094_),
    .Z(_0034_));
 MUX2_X1 _4533_ (.A(pwdata[1]),
    .B(\mem[15] [1]),
    .S(_1094_),
    .Z(_0035_));
 MUX2_X1 _4534_ (.A(pwdata[2]),
    .B(\mem[15] [2]),
    .S(_1094_),
    .Z(_0036_));
 MUX2_X1 _4535_ (.A(pwdata[3]),
    .B(\mem[15] [3]),
    .S(_1094_),
    .Z(_0037_));
 MUX2_X1 _4536_ (.A(pwdata[4]),
    .B(\mem[15] [4]),
    .S(_1094_),
    .Z(_0038_));
 MUX2_X1 _4537_ (.A(pwdata[5]),
    .B(\mem[15] [5]),
    .S(_1094_),
    .Z(_0039_));
 MUX2_X1 _4538_ (.A(pwdata[6]),
    .B(\mem[15] [6]),
    .S(_1094_),
    .Z(_0040_));
 MUX2_X1 _4539_ (.A(pwdata[7]),
    .B(\mem[15] [7]),
    .S(_1094_),
    .Z(_0041_));
 MUX2_X1 _4540_ (.A(pwdata[8]),
    .B(\mem[15] [8]),
    .S(_1094_),
    .Z(_0042_));
 MUX2_X1 _4541_ (.A(pwdata[9]),
    .B(\mem[15] [9]),
    .S(_1094_),
    .Z(_0043_));
 MUX2_X1 _4542_ (.A(pwdata[10]),
    .B(\mem[15] [10]),
    .S(_1094_),
    .Z(_0044_));
 MUX2_X1 _4543_ (.A(pwdata[11]),
    .B(\mem[15] [11]),
    .S(_1094_),
    .Z(_0045_));
 MUX2_X1 _4544_ (.A(pwdata[12]),
    .B(\mem[15] [12]),
    .S(_1094_),
    .Z(_0046_));
 MUX2_X1 _4545_ (.A(pwdata[13]),
    .B(\mem[15] [13]),
    .S(_1094_),
    .Z(_0047_));
 MUX2_X1 _4546_ (.A(pwdata[14]),
    .B(\mem[15] [14]),
    .S(_1094_),
    .Z(_0048_));
 MUX2_X1 _4547_ (.A(pwdata[15]),
    .B(\mem[15] [15]),
    .S(_1094_),
    .Z(_0049_));
 MUX2_X1 _4548_ (.A(pwdata[16]),
    .B(\mem[15] [16]),
    .S(_1094_),
    .Z(_0050_));
 MUX2_X1 _4549_ (.A(pwdata[17]),
    .B(\mem[15] [17]),
    .S(_1094_),
    .Z(_0051_));
 MUX2_X1 _4550_ (.A(pwdata[18]),
    .B(\mem[15] [18]),
    .S(_1094_),
    .Z(_0052_));
 MUX2_X1 _4551_ (.A(pwdata[19]),
    .B(\mem[15] [19]),
    .S(_1094_),
    .Z(_0053_));
 MUX2_X1 _4552_ (.A(pwdata[20]),
    .B(\mem[15] [20]),
    .S(_1094_),
    .Z(_0054_));
 MUX2_X1 _4553_ (.A(pwdata[21]),
    .B(\mem[15] [21]),
    .S(_1094_),
    .Z(_0055_));
 MUX2_X1 _4554_ (.A(pwdata[22]),
    .B(\mem[15] [22]),
    .S(_1094_),
    .Z(_0056_));
 MUX2_X1 _4555_ (.A(pwdata[23]),
    .B(\mem[15] [23]),
    .S(_1094_),
    .Z(_0057_));
 MUX2_X1 _4556_ (.A(pwdata[24]),
    .B(\mem[15] [24]),
    .S(_1094_),
    .Z(_0058_));
 MUX2_X1 _4557_ (.A(pwdata[25]),
    .B(\mem[15] [25]),
    .S(_1094_),
    .Z(_0059_));
 MUX2_X1 _4558_ (.A(pwdata[26]),
    .B(\mem[15] [26]),
    .S(_1094_),
    .Z(_0060_));
 MUX2_X1 _4559_ (.A(pwdata[27]),
    .B(\mem[15] [27]),
    .S(_1094_),
    .Z(_0061_));
 MUX2_X1 _4560_ (.A(pwdata[28]),
    .B(\mem[15] [28]),
    .S(_1094_),
    .Z(_0062_));
 MUX2_X1 _4561_ (.A(pwdata[29]),
    .B(\mem[15] [29]),
    .S(_1094_),
    .Z(_0063_));
 MUX2_X1 _4562_ (.A(pwdata[30]),
    .B(\mem[15] [30]),
    .S(_1094_),
    .Z(_0064_));
 MUX2_X1 _4563_ (.A(pwdata[31]),
    .B(\mem[15] [31]),
    .S(_1094_),
    .Z(_0065_));
 NOR4_X1 _4564_ (.A1(_1070_),
    .A2(paddr[2]),
    .A3(_1072_),
    .A4(paddr[0]),
    .ZN(_1095_));
 AND2_X2 _4565_ (.A1(paddr[4]),
    .A2(_1095_),
    .ZN(_1096_));
 NAND2_X4 _4566_ (.A1(net2),
    .A2(_1096_),
    .ZN(_1097_));
 MUX2_X1 _4567_ (.A(pwdata[0]),
    .B(\mem[26] [0]),
    .S(_1097_),
    .Z(_0066_));
 MUX2_X1 _4568_ (.A(pwdata[1]),
    .B(\mem[26] [1]),
    .S(_1097_),
    .Z(_0067_));
 MUX2_X1 _4569_ (.A(pwdata[2]),
    .B(\mem[26] [2]),
    .S(_1097_),
    .Z(_0068_));
 MUX2_X1 _4570_ (.A(pwdata[3]),
    .B(\mem[26] [3]),
    .S(_1097_),
    .Z(_0069_));
 MUX2_X1 _4571_ (.A(pwdata[4]),
    .B(\mem[26] [4]),
    .S(_1097_),
    .Z(_0070_));
 MUX2_X1 _4572_ (.A(pwdata[5]),
    .B(\mem[26] [5]),
    .S(_1097_),
    .Z(_0071_));
 MUX2_X1 _4573_ (.A(pwdata[6]),
    .B(\mem[26] [6]),
    .S(_1097_),
    .Z(_0072_));
 MUX2_X1 _4574_ (.A(pwdata[7]),
    .B(\mem[26] [7]),
    .S(_1097_),
    .Z(_0073_));
 MUX2_X1 _4575_ (.A(pwdata[8]),
    .B(\mem[26] [8]),
    .S(_1097_),
    .Z(_0074_));
 MUX2_X1 _4576_ (.A(pwdata[9]),
    .B(\mem[26] [9]),
    .S(_1097_),
    .Z(_0075_));
 MUX2_X1 _4577_ (.A(pwdata[10]),
    .B(\mem[26] [10]),
    .S(_1097_),
    .Z(_0076_));
 MUX2_X1 _4578_ (.A(pwdata[11]),
    .B(\mem[26] [11]),
    .S(_1097_),
    .Z(_0077_));
 MUX2_X1 _4579_ (.A(pwdata[12]),
    .B(\mem[26] [12]),
    .S(_1097_),
    .Z(_0078_));
 MUX2_X1 _4580_ (.A(pwdata[13]),
    .B(\mem[26] [13]),
    .S(_1097_),
    .Z(_0079_));
 MUX2_X1 _4581_ (.A(pwdata[14]),
    .B(\mem[26] [14]),
    .S(_1097_),
    .Z(_0080_));
 MUX2_X1 _4582_ (.A(pwdata[15]),
    .B(\mem[26] [15]),
    .S(_1097_),
    .Z(_0081_));
 MUX2_X1 _4583_ (.A(pwdata[16]),
    .B(\mem[26] [16]),
    .S(_1097_),
    .Z(_0082_));
 MUX2_X1 _4584_ (.A(pwdata[17]),
    .B(\mem[26] [17]),
    .S(_1097_),
    .Z(_0083_));
 MUX2_X1 _4585_ (.A(pwdata[18]),
    .B(\mem[26] [18]),
    .S(_1097_),
    .Z(_0084_));
 MUX2_X1 _4586_ (.A(pwdata[19]),
    .B(\mem[26] [19]),
    .S(_1097_),
    .Z(_0085_));
 MUX2_X1 _4587_ (.A(pwdata[20]),
    .B(\mem[26] [20]),
    .S(_1097_),
    .Z(_0086_));
 MUX2_X1 _4588_ (.A(pwdata[21]),
    .B(\mem[26] [21]),
    .S(_1097_),
    .Z(_0087_));
 MUX2_X1 _4589_ (.A(pwdata[22]),
    .B(\mem[26] [22]),
    .S(_1097_),
    .Z(_0088_));
 MUX2_X1 _4590_ (.A(pwdata[23]),
    .B(\mem[26] [23]),
    .S(_1097_),
    .Z(_0089_));
 MUX2_X1 _4591_ (.A(pwdata[24]),
    .B(\mem[26] [24]),
    .S(_1097_),
    .Z(_0090_));
 MUX2_X1 _4592_ (.A(pwdata[25]),
    .B(\mem[26] [25]),
    .S(_1097_),
    .Z(_0091_));
 MUX2_X1 _4593_ (.A(pwdata[26]),
    .B(\mem[26] [26]),
    .S(_1097_),
    .Z(_0092_));
 MUX2_X1 _4594_ (.A(pwdata[27]),
    .B(\mem[26] [27]),
    .S(_1097_),
    .Z(_0093_));
 MUX2_X1 _4595_ (.A(pwdata[28]),
    .B(\mem[26] [28]),
    .S(_1097_),
    .Z(_0094_));
 MUX2_X1 _4596_ (.A(pwdata[29]),
    .B(\mem[26] [29]),
    .S(_1097_),
    .Z(_0095_));
 MUX2_X1 _4597_ (.A(pwdata[30]),
    .B(\mem[26] [30]),
    .S(_1097_),
    .Z(_0096_));
 MUX2_X1 _4598_ (.A(pwdata[31]),
    .B(\mem[26] [31]),
    .S(_1097_),
    .Z(_0097_));
 OR2_X2 _4599_ (.A1(paddr[3]),
    .A2(paddr[2]),
    .ZN(_1098_));
 NOR3_X4 _4600_ (.A1(_1069_),
    .A2(_1076_),
    .A3(_1098_),
    .ZN(_1099_));
 NAND2_X4 _4601_ (.A1(net2),
    .A2(net10),
    .ZN(_1100_));
 MUX2_X1 _4602_ (.A(pwdata[0]),
    .B(\mem[16] [0]),
    .S(_1100_),
    .Z(_0098_));
 MUX2_X1 _4603_ (.A(pwdata[1]),
    .B(\mem[16] [1]),
    .S(_1100_),
    .Z(_0099_));
 MUX2_X1 _4604_ (.A(pwdata[2]),
    .B(\mem[16] [2]),
    .S(_1100_),
    .Z(_0100_));
 MUX2_X1 _4605_ (.A(pwdata[3]),
    .B(\mem[16] [3]),
    .S(_1100_),
    .Z(_0101_));
 MUX2_X1 _4606_ (.A(pwdata[4]),
    .B(\mem[16] [4]),
    .S(_1100_),
    .Z(_0102_));
 MUX2_X1 _4607_ (.A(pwdata[5]),
    .B(\mem[16] [5]),
    .S(_1100_),
    .Z(_0103_));
 MUX2_X1 _4608_ (.A(pwdata[6]),
    .B(\mem[16] [6]),
    .S(_1100_),
    .Z(_0104_));
 MUX2_X1 _4609_ (.A(pwdata[7]),
    .B(\mem[16] [7]),
    .S(_1100_),
    .Z(_0105_));
 MUX2_X1 _4610_ (.A(pwdata[8]),
    .B(\mem[16] [8]),
    .S(_1100_),
    .Z(_0106_));
 MUX2_X1 _4611_ (.A(pwdata[9]),
    .B(\mem[16] [9]),
    .S(_1100_),
    .Z(_0107_));
 MUX2_X1 _4612_ (.A(pwdata[10]),
    .B(\mem[16] [10]),
    .S(_1100_),
    .Z(_0108_));
 MUX2_X1 _4613_ (.A(pwdata[11]),
    .B(\mem[16] [11]),
    .S(_1100_),
    .Z(_0109_));
 MUX2_X1 _4614_ (.A(pwdata[12]),
    .B(\mem[16] [12]),
    .S(_1100_),
    .Z(_0110_));
 MUX2_X1 _4615_ (.A(pwdata[13]),
    .B(\mem[16] [13]),
    .S(_1100_),
    .Z(_0111_));
 MUX2_X1 _4616_ (.A(pwdata[14]),
    .B(\mem[16] [14]),
    .S(_1100_),
    .Z(_0112_));
 MUX2_X1 _4617_ (.A(pwdata[15]),
    .B(\mem[16] [15]),
    .S(_1100_),
    .Z(_0113_));
 MUX2_X1 _4618_ (.A(pwdata[16]),
    .B(\mem[16] [16]),
    .S(_1100_),
    .Z(_0114_));
 MUX2_X1 _4619_ (.A(pwdata[17]),
    .B(\mem[16] [17]),
    .S(_1100_),
    .Z(_0115_));
 MUX2_X1 _4620_ (.A(pwdata[18]),
    .B(\mem[16] [18]),
    .S(_1100_),
    .Z(_0116_));
 MUX2_X1 _4621_ (.A(pwdata[19]),
    .B(\mem[16] [19]),
    .S(_1100_),
    .Z(_0117_));
 MUX2_X1 _4622_ (.A(pwdata[20]),
    .B(\mem[16] [20]),
    .S(_1100_),
    .Z(_0118_));
 MUX2_X1 _4623_ (.A(pwdata[21]),
    .B(\mem[16] [21]),
    .S(_1100_),
    .Z(_0119_));
 MUX2_X1 _4624_ (.A(pwdata[22]),
    .B(\mem[16] [22]),
    .S(_1100_),
    .Z(_0120_));
 MUX2_X1 _4625_ (.A(pwdata[23]),
    .B(\mem[16] [23]),
    .S(_1100_),
    .Z(_0121_));
 MUX2_X1 _4626_ (.A(pwdata[24]),
    .B(\mem[16] [24]),
    .S(_1100_),
    .Z(_0122_));
 MUX2_X1 _4627_ (.A(pwdata[25]),
    .B(\mem[16] [25]),
    .S(_1100_),
    .Z(_0123_));
 MUX2_X1 _4628_ (.A(pwdata[26]),
    .B(\mem[16] [26]),
    .S(_1100_),
    .Z(_0124_));
 MUX2_X1 _4629_ (.A(pwdata[27]),
    .B(\mem[16] [27]),
    .S(_1100_),
    .Z(_0125_));
 MUX2_X1 _4630_ (.A(pwdata[28]),
    .B(\mem[16] [28]),
    .S(_1100_),
    .Z(_0126_));
 MUX2_X1 _4631_ (.A(pwdata[29]),
    .B(\mem[16] [29]),
    .S(_1100_),
    .Z(_0127_));
 MUX2_X1 _4632_ (.A(pwdata[30]),
    .B(\mem[16] [30]),
    .S(_1100_),
    .Z(_0128_));
 MUX2_X1 _4633_ (.A(pwdata[31]),
    .B(\mem[16] [31]),
    .S(_1100_),
    .Z(_0129_));
 NOR3_X4 _4634_ (.A1(_1069_),
    .A2(_1075_),
    .A3(_1092_),
    .ZN(_1101_));
 NAND2_X4 _4635_ (.A1(net2),
    .A2(net7),
    .ZN(_1102_));
 MUX2_X1 _4636_ (.A(pwdata[0]),
    .B(\mem[31] [0]),
    .S(_1102_),
    .Z(_0130_));
 MUX2_X1 _4637_ (.A(pwdata[1]),
    .B(\mem[31] [1]),
    .S(_1102_),
    .Z(_0131_));
 MUX2_X1 _4638_ (.A(pwdata[2]),
    .B(\mem[31] [2]),
    .S(_1102_),
    .Z(_0132_));
 MUX2_X1 _4639_ (.A(pwdata[3]),
    .B(\mem[31] [3]),
    .S(_1102_),
    .Z(_0133_));
 MUX2_X1 _4640_ (.A(pwdata[4]),
    .B(\mem[31] [4]),
    .S(_1102_),
    .Z(_0134_));
 MUX2_X1 _4641_ (.A(pwdata[5]),
    .B(\mem[31] [5]),
    .S(_1102_),
    .Z(_0135_));
 MUX2_X1 _4642_ (.A(pwdata[6]),
    .B(\mem[31] [6]),
    .S(_1102_),
    .Z(_0136_));
 MUX2_X1 _4643_ (.A(pwdata[7]),
    .B(\mem[31] [7]),
    .S(_1102_),
    .Z(_0137_));
 MUX2_X1 _4644_ (.A(pwdata[8]),
    .B(\mem[31] [8]),
    .S(_1102_),
    .Z(_0138_));
 MUX2_X1 _4645_ (.A(pwdata[9]),
    .B(\mem[31] [9]),
    .S(_1102_),
    .Z(_0139_));
 MUX2_X1 _4646_ (.A(pwdata[10]),
    .B(\mem[31] [10]),
    .S(_1102_),
    .Z(_0140_));
 MUX2_X1 _4647_ (.A(pwdata[11]),
    .B(\mem[31] [11]),
    .S(_1102_),
    .Z(_0141_));
 MUX2_X1 _4648_ (.A(pwdata[12]),
    .B(\mem[31] [12]),
    .S(_1102_),
    .Z(_0142_));
 MUX2_X1 _4649_ (.A(pwdata[13]),
    .B(\mem[31] [13]),
    .S(_1102_),
    .Z(_0143_));
 MUX2_X1 _4650_ (.A(pwdata[14]),
    .B(\mem[31] [14]),
    .S(_1102_),
    .Z(_0144_));
 MUX2_X1 _4651_ (.A(pwdata[15]),
    .B(\mem[31] [15]),
    .S(_1102_),
    .Z(_0145_));
 MUX2_X1 _4652_ (.A(pwdata[16]),
    .B(\mem[31] [16]),
    .S(_1102_),
    .Z(_0146_));
 MUX2_X1 _4653_ (.A(pwdata[17]),
    .B(\mem[31] [17]),
    .S(_1102_),
    .Z(_0147_));
 DFF_X1 _4654_ (.D(_0002_),
    .CK(clknet_leaf_18_pclk),
    .Q(\mem[12] [0]),
    .QN(_2852_));
 DFF_X1 _4655_ (.D(_0003_),
    .CK(clknet_leaf_26_pclk),
    .Q(\mem[12] [1]),
    .QN(_2851_));
 DFF_X1 _4656_ (.D(_0004_),
    .CK(clknet_leaf_12_pclk),
    .Q(\mem[12] [2]),
    .QN(_2850_));
 DFF_X1 _4657_ (.D(_0005_),
    .CK(clknet_leaf_15_pclk),
    .Q(\mem[12] [3]),
    .QN(_2849_));
 DFF_X1 _4658_ (.D(_0006_),
    .CK(clknet_leaf_22_pclk),
    .Q(\mem[12] [4]),
    .QN(_2848_));
 DFF_X1 _4659_ (.D(_0007_),
    .CK(clknet_leaf_10_pclk),
    .Q(\mem[12] [5]),
    .QN(_2847_));
 DFF_X1 _4660_ (.D(_0008_),
    .CK(clknet_leaf_2_pclk),
    .Q(\mem[12] [6]),
    .QN(_2846_));
 DFF_X1 _4661_ (.D(_0009_),
    .CK(clknet_leaf_28_pclk),
    .Q(\mem[12] [7]),
    .QN(_2845_));
 DFF_X1 _4662_ (.D(_0010_),
    .CK(clknet_leaf_34_pclk),
    .Q(\mem[12] [8]),
    .QN(_2844_));
 DFF_X1 _4663_ (.D(_0011_),
    .CK(clknet_leaf_1_pclk),
    .Q(\mem[12] [9]),
    .QN(_2843_));
 DFF_X1 _4664_ (.D(_0012_),
    .CK(clknet_leaf_17_pclk),
    .Q(\mem[12] [10]),
    .QN(_2842_));
 DFF_X1 _4665_ (.D(_0013_),
    .CK(clknet_leaf_6_pclk),
    .Q(\mem[12] [11]),
    .QN(_2841_));
 DFF_X1 _4666_ (.D(_0014_),
    .CK(clknet_leaf_3_pclk),
    .Q(\mem[12] [12]),
    .QN(_2840_));
 DFF_X1 _4667_ (.D(_0015_),
    .CK(clknet_leaf_29_pclk),
    .Q(\mem[12] [13]),
    .QN(_2839_));
 DFF_X1 _4668_ (.D(_0016_),
    .CK(clknet_leaf_25_pclk),
    .Q(\mem[12] [14]),
    .QN(_2838_));
 DFF_X1 _4669_ (.D(_0017_),
    .CK(clknet_leaf_24_pclk),
    .Q(\mem[12] [15]),
    .QN(_2837_));
 DFF_X1 _4670_ (.D(_0018_),
    .CK(clknet_leaf_3_pclk),
    .Q(\mem[12] [16]),
    .QN(_2836_));
 DFF_X1 _4671_ (.D(_0019_),
    .CK(clknet_leaf_11_pclk),
    .Q(\mem[12] [17]),
    .QN(_2835_));
 DFF_X1 _4672_ (.D(_0020_),
    .CK(clknet_leaf_8_pclk),
    .Q(\mem[12] [18]),
    .QN(_2834_));
 DFF_X1 _4673_ (.D(_0021_),
    .CK(clknet_leaf_6_pclk),
    .Q(\mem[12] [19]),
    .QN(_2833_));
 DFF_X1 _4674_ (.D(_0022_),
    .CK(clknet_leaf_34_pclk),
    .Q(\mem[12] [20]),
    .QN(_2832_));
 DFF_X1 _4675_ (.D(_0023_),
    .CK(clknet_leaf_15_pclk),
    .Q(\mem[12] [21]),
    .QN(_2831_));
 DFF_X1 _4676_ (.D(_0024_),
    .CK(clknet_leaf_8_pclk),
    .Q(\mem[12] [22]),
    .QN(_2830_));
 DFF_X1 _4677_ (.D(_0025_),
    .CK(clknet_leaf_21_pclk),
    .Q(\mem[12] [23]),
    .QN(_2829_));
 DFF_X1 _4678_ (.D(_0026_),
    .CK(clknet_leaf_16_pclk),
    .Q(\mem[12] [24]),
    .QN(_2828_));
 DFF_X1 _4679_ (.D(_0027_),
    .CK(clknet_leaf_20_pclk),
    .Q(\mem[12] [25]),
    .QN(_2827_));
 DFF_X1 _4680_ (.D(_0028_),
    .CK(clknet_leaf_8_pclk),
    .Q(\mem[12] [26]),
    .QN(_2826_));
 DFF_X1 _4681_ (.D(_0029_),
    .CK(clknet_leaf_0_pclk),
    .Q(\mem[12] [27]),
    .QN(_2825_));
 DFF_X1 _4682_ (.D(_0030_),
    .CK(clknet_leaf_29_pclk),
    .Q(\mem[12] [28]),
    .QN(_2824_));
 DFF_X1 _4683_ (.D(_0031_),
    .CK(clknet_leaf_32_pclk),
    .Q(\mem[12] [29]),
    .QN(_2823_));
 DFF_X1 _4684_ (.D(_0032_),
    .CK(clknet_leaf_19_pclk),
    .Q(\mem[12] [30]),
    .QN(_2822_));
 DFF_X1 _4685_ (.D(_0033_),
    .CK(clknet_leaf_28_pclk),
    .Q(\mem[12] [31]),
    .QN(_2853_));
 DFFR_X1 _4686_ (.D(_2855_[0]),
    .RN(prst_n),
    .CK(clknet_leaf_18_pclk),
    .Q(pready),
    .QN(_2821_));
 DFF_X1 _4687_ (.D(_0034_),
    .CK(clknet_leaf_18_pclk),
    .Q(\mem[15] [0]),
    .QN(_2820_));
 DFF_X1 _4688_ (.D(_0035_),
    .CK(clknet_leaf_27_pclk),
    .Q(\mem[15] [1]),
    .QN(_2819_));
 DFF_X1 _4689_ (.D(_0036_),
    .CK(clknet_leaf_30_pclk),
    .Q(\mem[15] [2]),
    .QN(_2818_));
 DFF_X1 _4690_ (.D(_0037_),
    .CK(clknet_leaf_14_pclk),
    .Q(\mem[15] [3]),
    .QN(_2817_));
 DFF_X1 _4691_ (.D(_0038_),
    .CK(clknet_leaf_23_pclk),
    .Q(\mem[15] [4]),
    .QN(_2816_));
 DFF_X1 _4692_ (.D(_0039_),
    .CK(clknet_leaf_10_pclk),
    .Q(\mem[15] [5]),
    .QN(_2815_));
 DFF_X1 _4693_ (.D(_0040_),
    .CK(clknet_leaf_1_pclk),
    .Q(\mem[15] [6]),
    .QN(_2814_));
 DFF_X1 _4694_ (.D(_0041_),
    .CK(clknet_leaf_28_pclk),
    .Q(\mem[15] [7]),
    .QN(_2813_));
 DFF_X1 _4695_ (.D(_0042_),
    .CK(clknet_leaf_34_pclk),
    .Q(\mem[15] [8]),
    .QN(_2812_));
 DFF_X1 _4696_ (.D(_0043_),
    .CK(clknet_leaf_5_pclk),
    .Q(\mem[15] [9]),
    .QN(_2811_));
 DFF_X1 _4697_ (.D(_0044_),
    .CK(clknet_leaf_18_pclk),
    .Q(\mem[15] [10]),
    .QN(_2810_));
 DFF_X1 _4698_ (.D(_0045_),
    .CK(clknet_leaf_4_pclk),
    .Q(\mem[15] [11]),
    .QN(_2809_));
 DFF_X1 _4699_ (.D(_0046_),
    .CK(clknet_leaf_2_pclk),
    .Q(\mem[15] [12]),
    .QN(_2808_));
 DFF_X1 _4700_ (.D(_0047_),
    .CK(clknet_leaf_29_pclk),
    .Q(\mem[15] [13]),
    .QN(_2807_));
 DFF_X1 _4701_ (.D(_0048_),
    .CK(clknet_leaf_26_pclk),
    .Q(\mem[15] [14]),
    .QN(_2806_));
 DFF_X1 _4702_ (.D(_0049_),
    .CK(clknet_leaf_24_pclk),
    .Q(\mem[15] [15]),
    .QN(_2805_));
 DFF_X1 _4703_ (.D(_0050_),
    .CK(clknet_leaf_4_pclk),
    .Q(\mem[15] [16]),
    .QN(_2804_));
 DFF_X1 _4704_ (.D(_0051_),
    .CK(clknet_leaf_13_pclk),
    .Q(\mem[15] [17]),
    .QN(_2803_));
 DFF_X1 _4705_ (.D(_0052_),
    .CK(clknet_leaf_9_pclk),
    .Q(\mem[15] [18]),
    .QN(_2802_));
 DFF_X1 _4706_ (.D(_0053_),
    .CK(clknet_leaf_5_pclk),
    .Q(\mem[15] [19]),
    .QN(_2801_));
 DFF_X1 _4707_ (.D(_0054_),
    .CK(clknet_leaf_32_pclk),
    .Q(\mem[15] [20]),
    .QN(_2800_));
 DFF_X1 _4708_ (.D(_0055_),
    .CK(clknet_leaf_15_pclk),
    .Q(\mem[15] [21]),
    .QN(_2799_));
 DFF_X1 _4709_ (.D(_0056_),
    .CK(clknet_leaf_7_pclk),
    .Q(\mem[15] [22]),
    .QN(_2798_));
 DFF_X1 _4710_ (.D(_0057_),
    .CK(clknet_leaf_30_pclk),
    .Q(\mem[15] [23]),
    .QN(_2797_));
 DFF_X1 _4711_ (.D(_0058_),
    .CK(clknet_leaf_16_pclk),
    .Q(\mem[15] [24]),
    .QN(_2796_));
 DFF_X1 _4712_ (.D(_0059_),
    .CK(clknet_leaf_20_pclk),
    .Q(\mem[15] [25]),
    .QN(_2795_));
 DFF_X1 _4713_ (.D(_0060_),
    .CK(clknet_leaf_8_pclk),
    .Q(\mem[15] [26]),
    .QN(_2794_));
 DFF_X1 _4714_ (.D(_0061_),
    .CK(clknet_leaf_0_pclk),
    .Q(\mem[15] [27]),
    .QN(_2793_));
 DFF_X1 _4715_ (.D(_0062_),
    .CK(clknet_leaf_23_pclk),
    .Q(\mem[15] [28]),
    .QN(_2792_));
 DFF_X1 _4716_ (.D(_0063_),
    .CK(clknet_leaf_32_pclk),
    .Q(\mem[15] [29]),
    .QN(_2791_));
 DFF_X1 _4717_ (.D(_0064_),
    .CK(clknet_leaf_18_pclk),
    .Q(\mem[15] [30]),
    .QN(_2790_));
 DFF_X1 _4718_ (.D(_0065_),
    .CK(clknet_leaf_32_pclk),
    .Q(\mem[15] [31]),
    .QN(_2789_));
 DFF_X1 _4719_ (.D(_0066_),
    .CK(clknet_leaf_19_pclk),
    .Q(\mem[26] [0]),
    .QN(_2788_));
 DFF_X1 _4720_ (.D(_0067_),
    .CK(clknet_leaf_26_pclk),
    .Q(\mem[26] [1]),
    .QN(_2787_));
 DFF_X1 _4721_ (.D(_0068_),
    .CK(clknet_leaf_3_pclk),
    .Q(\mem[26] [2]),
    .QN(_2786_));
 DFF_X1 _4722_ (.D(_0069_),
    .CK(clknet_leaf_14_pclk),
    .Q(\mem[26] [3]),
    .QN(_2785_));
 DFF_X1 _4723_ (.D(_0070_),
    .CK(clknet_leaf_23_pclk),
    .Q(\mem[26] [4]),
    .QN(_2784_));
 DFF_X1 _4724_ (.D(_0071_),
    .CK(clknet_leaf_10_pclk),
    .Q(\mem[26] [5]),
    .QN(_2783_));
 DFF_X1 _4725_ (.D(_0072_),
    .CK(clknet_leaf_1_pclk),
    .Q(\mem[26] [6]),
    .QN(_2782_));
 DFF_X1 _4726_ (.D(_0073_),
    .CK(clknet_leaf_28_pclk),
    .Q(\mem[26] [7]),
    .QN(_2781_));
 DFF_X1 _4727_ (.D(_0074_),
    .CK(clknet_leaf_33_pclk),
    .Q(\mem[26] [8]),
    .QN(_2780_));
 DFF_X1 _4728_ (.D(_0075_),
    .CK(clknet_leaf_2_pclk),
    .Q(\mem[26] [9]),
    .QN(_2779_));
 DFF_X1 _4729_ (.D(_0076_),
    .CK(clknet_leaf_16_pclk),
    .Q(\mem[26] [10]),
    .QN(_2778_));
 DFF_X1 _4730_ (.D(_0077_),
    .CK(clknet_leaf_6_pclk),
    .Q(\mem[26] [11]),
    .QN(_2777_));
 DFF_X1 _4731_ (.D(_0078_),
    .CK(clknet_leaf_31_pclk),
    .Q(\mem[26] [12]),
    .QN(_2776_));
 DFF_X1 _4732_ (.D(_0079_),
    .CK(clknet_leaf_22_pclk),
    .Q(\mem[26] [13]),
    .QN(_2775_));
 DFF_X1 _4733_ (.D(_0080_),
    .CK(clknet_leaf_24_pclk),
    .Q(\mem[26] [14]),
    .QN(_2774_));
 DFF_X1 _4734_ (.D(_0081_),
    .CK(clknet_leaf_24_pclk),
    .Q(\mem[26] [15]),
    .QN(_2773_));
 DFF_X1 _4735_ (.D(_0082_),
    .CK(clknet_leaf_11_pclk),
    .Q(\mem[26] [16]),
    .QN(_2772_));
 DFF_X1 _4736_ (.D(_0083_),
    .CK(clknet_leaf_13_pclk),
    .Q(\mem[26] [17]),
    .QN(_2771_));
 DFF_X1 _4737_ (.D(_0084_),
    .CK(clknet_leaf_9_pclk),
    .Q(\mem[26] [18]),
    .QN(_2770_));
 DFF_X1 _4738_ (.D(_0085_),
    .CK(clknet_leaf_6_pclk),
    .Q(\mem[26] [19]),
    .QN(_2769_));
 DFF_X1 _4739_ (.D(_0086_),
    .CK(clknet_leaf_33_pclk),
    .Q(\mem[26] [20]),
    .QN(_2768_));
 DFF_X1 _4740_ (.D(_0087_),
    .CK(clknet_leaf_20_pclk),
    .Q(\mem[26] [21]),
    .QN(_2767_));
 DFF_X1 _4741_ (.D(_0088_),
    .CK(clknet_leaf_8_pclk),
    .Q(\mem[26] [22]),
    .QN(_2766_));
 DFF_X1 _4742_ (.D(_0089_),
    .CK(clknet_leaf_30_pclk),
    .Q(\mem[26] [23]),
    .QN(_2765_));
 DFF_X1 _4743_ (.D(_0090_),
    .CK(clknet_leaf_16_pclk),
    .Q(\mem[26] [24]),
    .QN(_2764_));
 DFF_X1 _4744_ (.D(_0091_),
    .CK(clknet_leaf_21_pclk),
    .Q(\mem[26] [25]),
    .QN(_2763_));
 DFF_X1 _4745_ (.D(_0092_),
    .CK(clknet_leaf_9_pclk),
    .Q(\mem[26] [26]),
    .QN(_2762_));
 DFF_X1 _4746_ (.D(_0093_),
    .CK(clknet_leaf_0_pclk),
    .Q(\mem[26] [27]),
    .QN(_2761_));
 DFF_X1 _4747_ (.D(_0094_),
    .CK(clknet_leaf_24_pclk),
    .Q(\mem[26] [28]),
    .QN(_2760_));
 DFF_X1 _4748_ (.D(_0095_),
    .CK(clknet_leaf_31_pclk),
    .Q(\mem[26] [29]),
    .QN(_2759_));
 DFF_X1 _4749_ (.D(_0096_),
    .CK(clknet_leaf_23_pclk),
    .Q(\mem[26] [30]),
    .QN(_2758_));
 DFF_X1 _4750_ (.D(_0097_),
    .CK(clknet_leaf_28_pclk),
    .Q(\mem[26] [31]),
    .QN(_2757_));
 DFF_X1 _4751_ (.D(_0098_),
    .CK(clknet_leaf_18_pclk),
    .Q(\mem[16] [0]),
    .QN(_2756_));
 DFF_X1 _4752_ (.D(_0099_),
    .CK(clknet_leaf_27_pclk),
    .Q(\mem[16] [1]),
    .QN(_2755_));
 DFF_X1 _4753_ (.D(_0100_),
    .CK(clknet_leaf_3_pclk),
    .Q(\mem[16] [2]),
    .QN(_2754_));
 DFF_X1 _4754_ (.D(_0101_),
    .CK(clknet_leaf_13_pclk),
    .Q(\mem[16] [3]),
    .QN(_2753_));
 DFF_X1 _4755_ (.D(_0102_),
    .CK(clknet_leaf_23_pclk),
    .Q(\mem[16] [4]),
    .QN(_2752_));
 DFF_X1 _4756_ (.D(_0103_),
    .CK(clknet_leaf_10_pclk),
    .Q(\mem[16] [5]),
    .QN(_2751_));
 DFF_X1 _4757_ (.D(_0104_),
    .CK(clknet_leaf_2_pclk),
    .Q(\mem[16] [6]),
    .QN(_2750_));
 DFF_X1 _4758_ (.D(_0105_),
    .CK(clknet_leaf_27_pclk),
    .Q(\mem[16] [7]),
    .QN(_2749_));
 DFF_X1 _4759_ (.D(_0106_),
    .CK(clknet_leaf_34_pclk),
    .Q(\mem[16] [8]),
    .QN(_2748_));
 DFF_X1 _4760_ (.D(_0107_),
    .CK(clknet_leaf_5_pclk),
    .Q(\mem[16] [9]),
    .QN(_2747_));
 DFF_X1 _4761_ (.D(_0108_),
    .CK(clknet_leaf_18_pclk),
    .Q(\mem[16] [10]),
    .QN(_2746_));
 DFF_X1 _4762_ (.D(_0109_),
    .CK(clknet_leaf_5_pclk),
    .Q(\mem[16] [11]),
    .QN(_2745_));
 DFF_X1 _4763_ (.D(_0110_),
    .CK(clknet_leaf_31_pclk),
    .Q(\mem[16] [12]),
    .QN(_2744_));
 DFF_X1 _4764_ (.D(_0111_),
    .CK(clknet_leaf_29_pclk),
    .Q(\mem[16] [13]),
    .QN(_2743_));
 DFF_X1 _4765_ (.D(_0112_),
    .CK(clknet_leaf_25_pclk),
    .Q(\mem[16] [14]),
    .QN(_2742_));
 DFF_X1 _4766_ (.D(_0113_),
    .CK(clknet_leaf_24_pclk),
    .Q(\mem[16] [15]),
    .QN(_2741_));
 DFF_X1 _4767_ (.D(_0114_),
    .CK(clknet_leaf_11_pclk),
    .Q(\mem[16] [16]),
    .QN(_2740_));
 DFF_X1 _4768_ (.D(_0115_),
    .CK(clknet_leaf_12_pclk),
    .Q(\mem[16] [17]),
    .QN(_2739_));
 DFF_X1 _4769_ (.D(_0116_),
    .CK(clknet_leaf_11_pclk),
    .Q(\mem[16] [18]),
    .QN(_2738_));
 DFF_X1 _4770_ (.D(_0117_),
    .CK(clknet_leaf_6_pclk),
    .Q(\mem[16] [19]),
    .QN(_2737_));
 DFF_X1 _4771_ (.D(_0118_),
    .CK(clknet_leaf_33_pclk),
    .Q(\mem[16] [20]),
    .QN(_2736_));
 DFF_X1 _4772_ (.D(_0119_),
    .CK(clknet_leaf_15_pclk),
    .Q(\mem[16] [21]),
    .QN(_2735_));
 DFF_X1 _4773_ (.D(_0120_),
    .CK(clknet_leaf_8_pclk),
    .Q(\mem[16] [22]),
    .QN(_2734_));
 DFF_X1 _4774_ (.D(_0121_),
    .CK(clknet_leaf_30_pclk),
    .Q(\mem[16] [23]),
    .QN(_2733_));
 DFF_X1 _4775_ (.D(_0122_),
    .CK(clknet_leaf_17_pclk),
    .Q(\mem[16] [24]),
    .QN(_2732_));
 DFF_X1 _4776_ (.D(_0123_),
    .CK(clknet_leaf_21_pclk),
    .Q(\mem[16] [25]),
    .QN(_2731_));
 DFF_X1 _4777_ (.D(_0124_),
    .CK(clknet_leaf_9_pclk),
    .Q(\mem[16] [26]),
    .QN(_2730_));
 DFF_X1 _4778_ (.D(_0125_),
    .CK(clknet_leaf_0_pclk),
    .Q(\mem[16] [27]),
    .QN(_2729_));
 DFF_X1 _4779_ (.D(_0126_),
    .CK(clknet_leaf_23_pclk),
    .Q(\mem[16] [28]),
    .QN(_2728_));
 DFF_X1 _4780_ (.D(_0127_),
    .CK(clknet_leaf_33_pclk),
    .Q(\mem[16] [29]),
    .QN(_2727_));
 DFF_X1 _4781_ (.D(_0128_),
    .CK(clknet_leaf_19_pclk),
    .Q(\mem[16] [30]),
    .QN(_2726_));
 DFF_X1 _4782_ (.D(_0129_),
    .CK(clknet_leaf_31_pclk),
    .Q(\mem[16] [31]),
    .QN(_2725_));
 DFF_X1 _4783_ (.D(_0130_),
    .CK(clknet_leaf_20_pclk),
    .Q(\mem[31] [0]),
    .QN(_2724_));
 DFF_X1 _4784_ (.D(_0131_),
    .CK(clknet_leaf_26_pclk),
    .Q(\mem[31] [1]),
    .QN(_2723_));
 DFF_X1 _4785_ (.D(_0132_),
    .CK(clknet_leaf_3_pclk),
    .Q(\mem[31] [2]),
    .QN(_2722_));
 DFF_X1 _4786_ (.D(_0133_),
    .CK(clknet_leaf_15_pclk),
    .Q(\mem[31] [3]),
    .QN(_2721_));
 DFF_X1 _4787_ (.D(_0134_),
    .CK(clknet_leaf_21_pclk),
    .Q(\mem[31] [4]),
    .QN(_2720_));
 DFF_X1 _4788_ (.D(_0135_),
    .CK(clknet_leaf_10_pclk),
    .Q(\mem[31] [5]),
    .QN(_2719_));
 DFF_X1 _4789_ (.D(_0136_),
    .CK(clknet_leaf_2_pclk),
    .Q(\mem[31] [6]),
    .QN(_2718_));
 DFF_X1 _4790_ (.D(_0137_),
    .CK(clknet_leaf_28_pclk),
    .Q(\mem[31] [7]),
    .QN(_2717_));
 DFF_X1 _4791_ (.D(_0138_),
    .CK(clknet_leaf_35_pclk),
    .Q(\mem[31] [8]),
    .QN(_2716_));
 DFF_X1 _4792_ (.D(_0139_),
    .CK(clknet_leaf_5_pclk),
    .Q(\mem[31] [9]),
    .QN(_2715_));
 DFF_X1 _4793_ (.D(_0140_),
    .CK(clknet_leaf_17_pclk),
    .Q(\mem[31] [10]),
    .QN(_2714_));
 DFF_X1 _4794_ (.D(_0141_),
    .CK(clknet_leaf_4_pclk),
    .Q(\mem[31] [11]),
    .QN(_2713_));
 DFF_X1 _4795_ (.D(_0142_),
    .CK(clknet_leaf_3_pclk),
    .Q(\mem[31] [12]),
    .QN(_2712_));
 DFF_X1 _4796_ (.D(_0143_),
    .CK(clknet_leaf_22_pclk),
    .Q(\mem[31] [13]),
    .QN(_2711_));
 DFF_X1 _4797_ (.D(_0144_),
    .CK(clknet_leaf_26_pclk),
    .Q(\mem[31] [14]),
    .QN(_2710_));
 DFF_X1 _4798_ (.D(_0145_),
    .CK(clknet_leaf_24_pclk),
    .Q(\mem[31] [15]),
    .QN(_2709_));
 DFF_X1 _4799_ (.D(_0146_),
    .CK(clknet_leaf_11_pclk),
    .Q(\mem[31] [16]),
    .QN(_2708_));
 DFF_X1 _4800_ (.D(_0147_),
    .CK(clknet_leaf_14_pclk),
    .Q(\mem[31] [17]),
    .QN(_2707_));
 DFF_X1 _4801_ (.D(_0148_),
    .CK(clknet_leaf_9_pclk),
    .Q(\mem[31] [18]),
    .QN(_2706_));
 DFF_X1 _4802_ (.D(_0149_),
    .CK(clknet_leaf_6_pclk),
    .Q(\mem[31] [19]),
    .QN(_2705_));
 DFF_X1 _4803_ (.D(_0150_),
    .CK(clknet_leaf_33_pclk),
    .Q(\mem[31] [20]),
    .QN(_2704_));
 DFF_X1 _4804_ (.D(_0151_),
    .CK(clknet_leaf_13_pclk),
    .Q(\mem[31] [21]),
    .QN(_2703_));
 DFF_X1 _4805_ (.D(_0152_),
    .CK(clknet_leaf_8_pclk),
    .Q(\mem[31] [22]),
    .QN(_2702_));
 DFF_X1 _4806_ (.D(_0153_),
    .CK(clknet_leaf_3_pclk),
    .Q(\mem[31] [23]),
    .QN(_2701_));
 DFF_X1 _4807_ (.D(_0154_),
    .CK(clknet_leaf_16_pclk),
    .Q(\mem[31] [24]),
    .QN(_2700_));
 DFF_X1 _4808_ (.D(_0155_),
    .CK(clknet_leaf_20_pclk),
    .Q(\mem[31] [25]),
    .QN(_2699_));
 DFF_X1 _4809_ (.D(_0156_),
    .CK(clknet_leaf_8_pclk),
    .Q(\mem[31] [26]),
    .QN(_2698_));
 DFF_X1 _4810_ (.D(_0157_),
    .CK(clknet_leaf_0_pclk),
    .Q(\mem[31] [27]),
    .QN(_2697_));
 DFF_X1 _4811_ (.D(_0158_),
    .CK(clknet_leaf_22_pclk),
    .Q(\mem[31] [28]),
    .QN(_2696_));
 DFF_X1 _4812_ (.D(_0159_),
    .CK(clknet_leaf_32_pclk),
    .Q(\mem[31] [29]),
    .QN(_2695_));
 DFF_X1 _4813_ (.D(_0160_),
    .CK(clknet_leaf_22_pclk),
    .Q(\mem[31] [30]),
    .QN(_2694_));
 DFF_X1 _4814_ (.D(_0161_),
    .CK(clknet_leaf_28_pclk),
    .Q(\mem[31] [31]),
    .QN(_2693_));
 DFF_X1 _4815_ (.D(_0162_),
    .CK(clknet_leaf_18_pclk),
    .Q(\mem[17] [0]),
    .QN(_2692_));
 DFF_X1 _4816_ (.D(_0163_),
    .CK(clknet_leaf_27_pclk),
    .Q(\mem[17] [1]),
    .QN(_2691_));
 DFF_X1 _4817_ (.D(_0164_),
    .CK(clknet_leaf_3_pclk),
    .Q(\mem[17] [2]),
    .QN(_2690_));
 DFF_X1 _4818_ (.D(_0165_),
    .CK(clknet_leaf_13_pclk),
    .Q(\mem[17] [3]),
    .QN(_2689_));
 DFF_X1 _4819_ (.D(_0166_),
    .CK(clknet_leaf_23_pclk),
    .Q(\mem[17] [4]),
    .QN(_2688_));
 DFF_X1 _4820_ (.D(_0167_),
    .CK(clknet_leaf_10_pclk),
    .Q(\mem[17] [5]),
    .QN(_2687_));
 DFF_X1 _4821_ (.D(_0168_),
    .CK(clknet_leaf_2_pclk),
    .Q(\mem[17] [6]),
    .QN(_2686_));
 DFF_X1 _4822_ (.D(_0169_),
    .CK(clknet_leaf_27_pclk),
    .Q(\mem[17] [7]),
    .QN(_2685_));
 DFF_X1 _4823_ (.D(_0170_),
    .CK(clknet_leaf_34_pclk),
    .Q(\mem[17] [8]),
    .QN(_2684_));
 DFF_X1 _4824_ (.D(_0171_),
    .CK(clknet_leaf_5_pclk),
    .Q(\mem[17] [9]),
    .QN(_2683_));
 DFF_X1 _4825_ (.D(_0172_),
    .CK(clknet_leaf_17_pclk),
    .Q(\mem[17] [10]),
    .QN(_2682_));
 DFF_X1 _4826_ (.D(_0173_),
    .CK(clknet_leaf_6_pclk),
    .Q(\mem[17] [11]),
    .QN(_2681_));
 DFF_X1 _4827_ (.D(_0174_),
    .CK(clknet_leaf_30_pclk),
    .Q(\mem[17] [12]),
    .QN(_2680_));
 DFF_X1 _4828_ (.D(_0175_),
    .CK(clknet_leaf_21_pclk),
    .Q(\mem[17] [13]),
    .QN(_2679_));
 DFF_X1 _4829_ (.D(_0176_),
    .CK(clknet_leaf_25_pclk),
    .Q(\mem[17] [14]),
    .QN(_2678_));
 DFF_X1 _4830_ (.D(_0177_),
    .CK(clknet_leaf_24_pclk),
    .Q(\mem[17] [15]),
    .QN(_2677_));
 DFF_X1 _4831_ (.D(_0178_),
    .CK(clknet_leaf_4_pclk),
    .Q(\mem[17] [16]),
    .QN(_2676_));
 DFF_X1 _4832_ (.D(_0179_),
    .CK(clknet_leaf_12_pclk),
    .Q(\mem[17] [17]),
    .QN(_2675_));
 DFF_X1 _4833_ (.D(_0180_),
    .CK(clknet_leaf_11_pclk),
    .Q(\mem[17] [18]),
    .QN(_2674_));
 DFF_X1 _4834_ (.D(_0181_),
    .CK(clknet_leaf_5_pclk),
    .Q(\mem[17] [19]),
    .QN(_2673_));
 DFF_X1 _4835_ (.D(_0182_),
    .CK(clknet_leaf_34_pclk),
    .Q(\mem[17] [20]),
    .QN(_2672_));
 DFF_X1 _4836_ (.D(_0183_),
    .CK(clknet_leaf_15_pclk),
    .Q(\mem[17] [21]),
    .QN(_2671_));
 DFF_X1 _4837_ (.D(_0184_),
    .CK(clknet_leaf_7_pclk),
    .Q(\mem[17] [22]),
    .QN(_2670_));
 DFF_X1 _4838_ (.D(_0185_),
    .CK(clknet_leaf_30_pclk),
    .Q(\mem[17] [23]),
    .QN(_2669_));
 DFF_X1 _4839_ (.D(_0186_),
    .CK(clknet_leaf_17_pclk),
    .Q(\mem[17] [24]),
    .QN(_2668_));
 DFF_X1 _4840_ (.D(_0187_),
    .CK(clknet_leaf_20_pclk),
    .Q(\mem[17] [25]),
    .QN(_2667_));
 DFF_X1 _4841_ (.D(_0188_),
    .CK(clknet_leaf_7_pclk),
    .Q(\mem[17] [26]),
    .QN(_2666_));
 DFF_X1 _4842_ (.D(_0189_),
    .CK(clknet_leaf_1_pclk),
    .Q(\mem[17] [27]),
    .QN(_2665_));
 DFF_X1 _4843_ (.D(_0190_),
    .CK(clknet_leaf_28_pclk),
    .Q(\mem[17] [28]),
    .QN(_2664_));
 DFF_X1 _4844_ (.D(_0191_),
    .CK(clknet_leaf_32_pclk),
    .Q(\mem[17] [29]),
    .QN(_2663_));
 DFF_X1 _4845_ (.D(_0192_),
    .CK(clknet_leaf_19_pclk),
    .Q(\mem[17] [30]),
    .QN(_2662_));
 DFF_X1 _4846_ (.D(_0193_),
    .CK(clknet_leaf_28_pclk),
    .Q(\mem[17] [31]),
    .QN(_2661_));
 DFF_X1 _4847_ (.D(_0194_),
    .CK(clknet_leaf_19_pclk),
    .Q(\mem[27] [0]),
    .QN(_2660_));
 DFF_X1 _4848_ (.D(_0195_),
    .CK(clknet_leaf_26_pclk),
    .Q(\mem[27] [1]),
    .QN(_2659_));
 DFF_X1 _4849_ (.D(_0196_),
    .CK(clknet_leaf_3_pclk),
    .Q(\mem[27] [2]),
    .QN(_2658_));
 DFF_X1 _4850_ (.D(_0197_),
    .CK(clknet_leaf_14_pclk),
    .Q(\mem[27] [3]),
    .QN(_2657_));
 DFF_X1 _4851_ (.D(_0198_),
    .CK(clknet_leaf_23_pclk),
    .Q(\mem[27] [4]),
    .QN(_2656_));
 DFF_X1 _4852_ (.D(_0199_),
    .CK(clknet_leaf_10_pclk),
    .Q(\mem[27] [5]),
    .QN(_2655_));
 DFF_X1 _4853_ (.D(_0200_),
    .CK(clknet_leaf_2_pclk),
    .Q(\mem[27] [6]),
    .QN(_2654_));
 DFF_X1 _4854_ (.D(_0201_),
    .CK(clknet_leaf_28_pclk),
    .Q(\mem[27] [7]),
    .QN(_2653_));
 DFF_X1 _4855_ (.D(_0202_),
    .CK(clknet_leaf_35_pclk),
    .Q(\mem[27] [8]),
    .QN(_2652_));
 DFF_X1 _4856_ (.D(_0203_),
    .CK(clknet_leaf_2_pclk),
    .Q(\mem[27] [9]),
    .QN(_2651_));
 DFF_X1 _4857_ (.D(_0204_),
    .CK(clknet_leaf_16_pclk),
    .Q(\mem[27] [10]),
    .QN(_2650_));
 DFF_X1 _4858_ (.D(_0205_),
    .CK(clknet_leaf_6_pclk),
    .Q(\mem[27] [11]),
    .QN(_2649_));
 DFF_X1 _4859_ (.D(_0206_),
    .CK(clknet_leaf_31_pclk),
    .Q(\mem[27] [12]),
    .QN(_2648_));
 DFF_X1 _4860_ (.D(_0207_),
    .CK(clknet_leaf_29_pclk),
    .Q(\mem[27] [13]),
    .QN(_2647_));
 DFF_X1 _4861_ (.D(_0208_),
    .CK(clknet_leaf_25_pclk),
    .Q(\mem[27] [14]),
    .QN(_2646_));
 DFF_X1 _4862_ (.D(_0209_),
    .CK(clknet_leaf_26_pclk),
    .Q(\mem[27] [15]),
    .QN(_2645_));
 DFF_X1 _4863_ (.D(_0210_),
    .CK(clknet_leaf_11_pclk),
    .Q(\mem[27] [16]),
    .QN(_2644_));
 DFF_X1 _4864_ (.D(_0211_),
    .CK(clknet_leaf_12_pclk),
    .Q(\mem[27] [17]),
    .QN(_2643_));
 DFF_X1 _4865_ (.D(_0212_),
    .CK(clknet_leaf_8_pclk),
    .Q(\mem[27] [18]),
    .QN(_2642_));
 DFF_X1 _4866_ (.D(_0213_),
    .CK(clknet_leaf_6_pclk),
    .Q(\mem[27] [19]),
    .QN(_2641_));
 DFF_X1 _4867_ (.D(_0214_),
    .CK(clknet_leaf_33_pclk),
    .Q(\mem[27] [20]),
    .QN(_2640_));
 DFF_X1 _4868_ (.D(_0215_),
    .CK(clknet_leaf_15_pclk),
    .Q(\mem[27] [21]),
    .QN(_2639_));
 DFF_X1 _4869_ (.D(_0216_),
    .CK(clknet_leaf_8_pclk),
    .Q(\mem[27] [22]),
    .QN(_2638_));
 DFF_X1 _4870_ (.D(_0217_),
    .CK(clknet_leaf_21_pclk),
    .Q(\mem[27] [23]),
    .QN(_2637_));
 DFF_X1 _4871_ (.D(_0218_),
    .CK(clknet_leaf_16_pclk),
    .Q(\mem[27] [24]),
    .QN(_2636_));
 DFF_X1 _4872_ (.D(_0219_),
    .CK(clknet_leaf_21_pclk),
    .Q(\mem[27] [25]),
    .QN(_2635_));
 DFF_X1 _4873_ (.D(_0220_),
    .CK(clknet_leaf_9_pclk),
    .Q(\mem[27] [26]),
    .QN(_2634_));
 DFF_X1 _4874_ (.D(_0221_),
    .CK(clknet_leaf_35_pclk),
    .Q(\mem[27] [27]),
    .QN(_2633_));
 DFF_X1 _4875_ (.D(_0222_),
    .CK(clknet_leaf_23_pclk),
    .Q(\mem[27] [28]),
    .QN(_2632_));
 DFF_X1 _4876_ (.D(_0223_),
    .CK(clknet_leaf_31_pclk),
    .Q(\mem[27] [29]),
    .QN(_2631_));
 DFF_X1 _4877_ (.D(_0224_),
    .CK(clknet_leaf_19_pclk),
    .Q(\mem[27] [30]),
    .QN(_2630_));
 DFF_X1 _4878_ (.D(_0225_),
    .CK(clknet_leaf_31_pclk),
    .Q(\mem[27] [31]),
    .QN(_2629_));
 DFF_X1 _4879_ (.D(_0226_),
    .CK(clknet_leaf_19_pclk),
    .Q(\mem[18] [0]),
    .QN(_2628_));
 DFF_X1 _4880_ (.D(_0227_),
    .CK(clknet_leaf_27_pclk),
    .Q(\mem[18] [1]),
    .QN(_2627_));
 DFF_X1 _4881_ (.D(_0228_),
    .CK(clknet_leaf_3_pclk),
    .Q(\mem[18] [2]),
    .QN(_2626_));
 DFF_X1 _4882_ (.D(_0229_),
    .CK(clknet_leaf_15_pclk),
    .Q(\mem[18] [3]),
    .QN(_2625_));
 DFF_X1 _4883_ (.D(_0230_),
    .CK(clknet_leaf_22_pclk),
    .Q(\mem[18] [4]),
    .QN(_2624_));
 DFF_X1 _4884_ (.D(_0231_),
    .CK(clknet_leaf_10_pclk),
    .Q(\mem[18] [5]),
    .QN(_2623_));
 DFF_X1 _4885_ (.D(_0232_),
    .CK(clknet_leaf_2_pclk),
    .Q(\mem[18] [6]),
    .QN(_2622_));
 DFF_X1 _4886_ (.D(_0233_),
    .CK(clknet_leaf_28_pclk),
    .Q(\mem[18] [7]),
    .QN(_2621_));
 DFF_X1 _4887_ (.D(_0234_),
    .CK(clknet_leaf_34_pclk),
    .Q(\mem[18] [8]),
    .QN(_2620_));
 DFF_X1 _4888_ (.D(_0235_),
    .CK(clknet_leaf_1_pclk),
    .Q(\mem[18] [9]),
    .QN(_2619_));
 DFF_X1 _4889_ (.D(_0236_),
    .CK(clknet_leaf_17_pclk),
    .Q(\mem[18] [10]),
    .QN(_2618_));
 DFF_X1 _4890_ (.D(_0237_),
    .CK(clknet_leaf_4_pclk),
    .Q(\mem[18] [11]),
    .QN(_2617_));
 DFF_X1 _4891_ (.D(_0238_),
    .CK(clknet_leaf_30_pclk),
    .Q(\mem[18] [12]),
    .QN(_2616_));
 DFF_X1 _4892_ (.D(_0239_),
    .CK(clknet_leaf_21_pclk),
    .Q(\mem[18] [13]),
    .QN(_2615_));
 DFF_X1 _4893_ (.D(_0240_),
    .CK(clknet_leaf_26_pclk),
    .Q(\mem[18] [14]),
    .QN(_2614_));
 DFF_X1 _4894_ (.D(_0241_),
    .CK(clknet_leaf_26_pclk),
    .Q(\mem[18] [15]),
    .QN(_2613_));
 DFF_X1 _4895_ (.D(_0242_),
    .CK(clknet_leaf_4_pclk),
    .Q(\mem[18] [16]),
    .QN(_2612_));
 DFF_X1 _4896_ (.D(_0243_),
    .CK(clknet_leaf_14_pclk),
    .Q(\mem[18] [17]),
    .QN(_2611_));
 DFF_X1 _4897_ (.D(_0244_),
    .CK(clknet_leaf_9_pclk),
    .Q(\mem[18] [18]),
    .QN(_2610_));
 DFF_X1 _4898_ (.D(_0245_),
    .CK(clknet_leaf_6_pclk),
    .Q(\mem[18] [19]),
    .QN(_2609_));
 DFF_X1 _4899_ (.D(_0246_),
    .CK(clknet_leaf_34_pclk),
    .Q(\mem[18] [20]),
    .QN(_2608_));
 DFF_X1 _4900_ (.D(_0247_),
    .CK(clknet_leaf_15_pclk),
    .Q(\mem[18] [21]),
    .QN(_2607_));
 DFF_X1 _4901_ (.D(_0248_),
    .CK(clknet_leaf_7_pclk),
    .Q(\mem[18] [22]),
    .QN(_2606_));
 DFF_X1 _4902_ (.D(_0249_),
    .CK(clknet_leaf_30_pclk),
    .Q(\mem[18] [23]),
    .QN(_2605_));
 DFF_X1 _4903_ (.D(_0250_),
    .CK(clknet_leaf_16_pclk),
    .Q(\mem[18] [24]),
    .QN(_2604_));
 DFF_X1 _4904_ (.D(_0251_),
    .CK(clknet_leaf_20_pclk),
    .Q(\mem[18] [25]),
    .QN(_2603_));
 DFF_X1 _4905_ (.D(_0252_),
    .CK(clknet_leaf_7_pclk),
    .Q(\mem[18] [26]),
    .QN(_2602_));
 DFF_X1 _4906_ (.D(_0253_),
    .CK(clknet_leaf_1_pclk),
    .Q(\mem[18] [27]),
    .QN(_2601_));
 DFF_X1 _4907_ (.D(_0254_),
    .CK(clknet_leaf_22_pclk),
    .Q(\mem[18] [28]),
    .QN(_2600_));
 DFF_X1 _4908_ (.D(_0255_),
    .CK(clknet_leaf_32_pclk),
    .Q(\mem[18] [29]),
    .QN(_2599_));
 DFF_X1 _4909_ (.D(_0256_),
    .CK(clknet_leaf_19_pclk),
    .Q(\mem[18] [30]),
    .QN(_2598_));
 DFF_X1 _4910_ (.D(_0257_),
    .CK(clknet_leaf_32_pclk),
    .Q(\mem[18] [31]),
    .QN(_2597_));
 DFF_X1 _4911_ (.D(_0258_),
    .CK(clknet_leaf_20_pclk),
    .Q(\mem[28] [0]),
    .QN(_2596_));
 DFF_X1 _4912_ (.D(_0259_),
    .CK(clknet_leaf_27_pclk),
    .Q(\mem[28] [1]),
    .QN(_2595_));
 DFF_X1 _4913_ (.D(_0260_),
    .CK(clknet_leaf_30_pclk),
    .Q(\mem[28] [2]),
    .QN(_2594_));
 DFF_X1 _4914_ (.D(_0261_),
    .CK(clknet_leaf_15_pclk),
    .Q(\mem[28] [3]),
    .QN(_2593_));
 DFF_X1 _4915_ (.D(_0262_),
    .CK(clknet_leaf_22_pclk),
    .Q(\mem[28] [4]),
    .QN(_2592_));
 DFF_X1 _4916_ (.D(_0263_),
    .CK(clknet_leaf_10_pclk),
    .Q(\mem[28] [5]),
    .QN(_2591_));
 DFF_X1 _4917_ (.D(_0264_),
    .CK(clknet_leaf_1_pclk),
    .Q(\mem[28] [6]),
    .QN(_2590_));
 DFF_X1 _4918_ (.D(_0265_),
    .CK(clknet_leaf_27_pclk),
    .Q(\mem[28] [7]),
    .QN(_2589_));
 DFF_X1 _4919_ (.D(_0266_),
    .CK(clknet_leaf_34_pclk),
    .Q(\mem[28] [8]),
    .QN(_2588_));
 DFF_X1 _4920_ (.D(_0267_),
    .CK(clknet_leaf_5_pclk),
    .Q(\mem[28] [9]),
    .QN(_2587_));
 DFF_X1 _4921_ (.D(_0268_),
    .CK(clknet_leaf_15_pclk),
    .Q(\mem[28] [10]),
    .QN(_2586_));
 DFF_X1 _4922_ (.D(_0269_),
    .CK(clknet_leaf_6_pclk),
    .Q(\mem[28] [11]),
    .QN(_2585_));
 DFF_X1 _4923_ (.D(_0270_),
    .CK(clknet_leaf_3_pclk),
    .Q(\mem[28] [12]),
    .QN(_2584_));
 DFF_X1 _4924_ (.D(_0271_),
    .CK(clknet_leaf_22_pclk),
    .Q(\mem[28] [13]),
    .QN(_2583_));
 DFF_X1 _4925_ (.D(_0272_),
    .CK(clknet_leaf_26_pclk),
    .Q(\mem[28] [14]),
    .QN(_2582_));
 DFF_X1 _4926_ (.D(_0273_),
    .CK(clknet_leaf_24_pclk),
    .Q(\mem[28] [15]),
    .QN(_2581_));
 DFF_X1 _4927_ (.D(_0274_),
    .CK(clknet_leaf_11_pclk),
    .Q(\mem[28] [16]),
    .QN(_2580_));
 DFF_X1 _4928_ (.D(_0275_),
    .CK(clknet_leaf_13_pclk),
    .Q(\mem[28] [17]),
    .QN(_2579_));
 DFF_X1 _4929_ (.D(_0276_),
    .CK(clknet_leaf_9_pclk),
    .Q(\mem[28] [18]),
    .QN(_2578_));
 DFF_X1 _4930_ (.D(_0277_),
    .CK(clknet_leaf_5_pclk),
    .Q(\mem[28] [19]),
    .QN(_2577_));
 DFF_X1 _4931_ (.D(_0278_),
    .CK(clknet_leaf_33_pclk),
    .Q(\mem[28] [20]),
    .QN(_2576_));
 DFF_X1 _4932_ (.D(_0279_),
    .CK(clknet_leaf_13_pclk),
    .Q(\mem[28] [21]),
    .QN(_2575_));
 DFF_X1 _4933_ (.D(_0280_),
    .CK(clknet_leaf_7_pclk),
    .Q(\mem[28] [22]),
    .QN(_2574_));
 DFF_X1 _4934_ (.D(_0281_),
    .CK(clknet_leaf_21_pclk),
    .Q(\mem[28] [23]),
    .QN(_2573_));
 DFF_X1 _4935_ (.D(_0282_),
    .CK(clknet_leaf_16_pclk),
    .Q(\mem[28] [24]),
    .QN(_2572_));
 DFF_X1 _4936_ (.D(_0283_),
    .CK(clknet_leaf_13_pclk),
    .Q(\mem[28] [25]),
    .QN(_2571_));
 DFF_X1 _4937_ (.D(_0284_),
    .CK(clknet_leaf_8_pclk),
    .Q(\mem[28] [26]),
    .QN(_2570_));
 DFF_X1 _4938_ (.D(_0285_),
    .CK(clknet_leaf_1_pclk),
    .Q(\mem[28] [27]),
    .QN(_2569_));
 DFF_X1 _4939_ (.D(_0286_),
    .CK(clknet_leaf_29_pclk),
    .Q(\mem[28] [28]),
    .QN(_2568_));
 DFF_X1 _4940_ (.D(_0287_),
    .CK(clknet_leaf_32_pclk),
    .Q(\mem[28] [29]),
    .QN(_2567_));
 DFF_X1 _4941_ (.D(_0288_),
    .CK(clknet_leaf_22_pclk),
    .Q(\mem[28] [30]),
    .QN(_2566_));
 DFF_X1 _4942_ (.D(_0289_),
    .CK(clknet_leaf_28_pclk),
    .Q(\mem[28] [31]),
    .QN(_2565_));
 DFF_X1 _4943_ (.D(_0290_),
    .CK(clknet_leaf_19_pclk),
    .Q(\mem[19] [0]),
    .QN(_2564_));
 DFF_X1 _4944_ (.D(_0291_),
    .CK(clknet_leaf_27_pclk),
    .Q(\mem[19] [1]),
    .QN(_2563_));
 DFF_X1 _4945_ (.D(_0292_),
    .CK(clknet_leaf_3_pclk),
    .Q(\mem[19] [2]),
    .QN(_2562_));
 DFF_X1 _4946_ (.D(_0293_),
    .CK(clknet_leaf_15_pclk),
    .Q(\mem[19] [3]),
    .QN(_2561_));
 DFF_X1 _4947_ (.D(_0294_),
    .CK(clknet_leaf_22_pclk),
    .Q(\mem[19] [4]),
    .QN(_2560_));
 DFF_X1 _4948_ (.D(_0295_),
    .CK(clknet_leaf_10_pclk),
    .Q(\mem[19] [5]),
    .QN(_2559_));
 DFF_X1 _4949_ (.D(_0296_),
    .CK(clknet_leaf_1_pclk),
    .Q(\mem[19] [6]),
    .QN(_2558_));
 DFF_X1 _4950_ (.D(_0297_),
    .CK(clknet_leaf_28_pclk),
    .Q(\mem[19] [7]),
    .QN(_2557_));
 DFF_X1 _4951_ (.D(_0298_),
    .CK(clknet_leaf_34_pclk),
    .Q(\mem[19] [8]),
    .QN(_2556_));
 DFF_X1 _4952_ (.D(_0299_),
    .CK(clknet_leaf_1_pclk),
    .Q(\mem[19] [9]),
    .QN(_2555_));
 DFF_X1 _4953_ (.D(_0300_),
    .CK(clknet_leaf_17_pclk),
    .Q(\mem[19] [10]),
    .QN(_2554_));
 DFF_X1 _4954_ (.D(_0301_),
    .CK(clknet_leaf_6_pclk),
    .Q(\mem[19] [11]),
    .QN(_2553_));
 DFF_X1 _4955_ (.D(_0302_),
    .CK(clknet_leaf_30_pclk),
    .Q(\mem[19] [12]),
    .QN(_2552_));
 DFF_X1 _4956_ (.D(_0303_),
    .CK(clknet_leaf_21_pclk),
    .Q(\mem[19] [13]),
    .QN(_2551_));
 DFF_X1 _4957_ (.D(_0304_),
    .CK(clknet_leaf_26_pclk),
    .Q(\mem[19] [14]),
    .QN(_2550_));
 DFF_X1 _4958_ (.D(_0305_),
    .CK(clknet_leaf_26_pclk),
    .Q(\mem[19] [15]),
    .QN(_2549_));
 DFF_X1 _4959_ (.D(_0306_),
    .CK(clknet_leaf_12_pclk),
    .Q(\mem[19] [16]),
    .QN(_2548_));
 DFF_X1 _4960_ (.D(_0307_),
    .CK(clknet_leaf_14_pclk),
    .Q(\mem[19] [17]),
    .QN(_2547_));
 DFF_X1 _4961_ (.D(_0308_),
    .CK(clknet_leaf_9_pclk),
    .Q(\mem[19] [18]),
    .QN(_2546_));
 DFF_X1 _4962_ (.D(_0309_),
    .CK(clknet_leaf_6_pclk),
    .Q(\mem[19] [19]),
    .QN(_2545_));
 DFF_X1 _4963_ (.D(_0310_),
    .CK(clknet_leaf_34_pclk),
    .Q(\mem[19] [20]),
    .QN(_2544_));
 DFF_X1 _4964_ (.D(_0311_),
    .CK(clknet_leaf_15_pclk),
    .Q(\mem[19] [21]),
    .QN(_2543_));
 DFF_X1 _4965_ (.D(_0312_),
    .CK(clknet_leaf_7_pclk),
    .Q(\mem[19] [22]),
    .QN(_2542_));
 DFF_X1 _4966_ (.D(_0313_),
    .CK(clknet_leaf_30_pclk),
    .Q(\mem[19] [23]),
    .QN(_2541_));
 DFF_X1 _4967_ (.D(_0314_),
    .CK(clknet_leaf_16_pclk),
    .Q(\mem[19] [24]),
    .QN(_2540_));
 DFF_X1 _4968_ (.D(_0315_),
    .CK(clknet_leaf_20_pclk),
    .Q(\mem[19] [25]),
    .QN(_2539_));
 DFF_X1 _4969_ (.D(_0316_),
    .CK(clknet_leaf_7_pclk),
    .Q(\mem[19] [26]),
    .QN(_2538_));
 DFF_X1 _4970_ (.D(_0317_),
    .CK(clknet_leaf_1_pclk),
    .Q(\mem[19] [27]),
    .QN(_2537_));
 DFF_X1 _4971_ (.D(_0318_),
    .CK(clknet_leaf_29_pclk),
    .Q(\mem[19] [28]),
    .QN(_2536_));
 DFF_X1 _4972_ (.D(_0319_),
    .CK(clknet_leaf_32_pclk),
    .Q(\mem[19] [29]),
    .QN(_2535_));
 DFF_X1 _4973_ (.D(_0320_),
    .CK(clknet_leaf_19_pclk),
    .Q(\mem[19] [30]),
    .QN(_2534_));
 DFF_X1 _4974_ (.D(_0321_),
    .CK(clknet_leaf_31_pclk),
    .Q(\mem[19] [31]),
    .QN(_2533_));
 DFF_X1 _4975_ (.D(_0322_),
    .CK(clknet_leaf_20_pclk),
    .Q(\mem[24] [0]),
    .QN(_2532_));
 DFF_X1 _4976_ (.D(_0323_),
    .CK(clknet_leaf_27_pclk),
    .Q(\mem[24] [1]),
    .QN(_2531_));
 DFF_X1 _4977_ (.D(_0324_),
    .CK(clknet_leaf_3_pclk),
    .Q(\mem[24] [2]),
    .QN(_2530_));
 DFF_X1 _4978_ (.D(_0325_),
    .CK(clknet_leaf_14_pclk),
    .Q(\mem[24] [3]),
    .QN(_2529_));
 DFF_X1 _4979_ (.D(_0326_),
    .CK(clknet_leaf_20_pclk),
    .Q(\mem[24] [4]),
    .QN(_2528_));
 DFF_X1 _4980_ (.D(_0327_),
    .CK(clknet_leaf_9_pclk),
    .Q(\mem[24] [5]),
    .QN(_2527_));
 DFF_X1 _4981_ (.D(_0328_),
    .CK(clknet_leaf_1_pclk),
    .Q(\mem[24] [6]),
    .QN(_2526_));
 DFF_X1 _4982_ (.D(_0329_),
    .CK(clknet_leaf_27_pclk),
    .Q(\mem[24] [7]),
    .QN(_2525_));
 DFF_X1 _4983_ (.D(_0330_),
    .CK(clknet_leaf_35_pclk),
    .Q(\mem[24] [8]),
    .QN(_2524_));
 DFF_X1 _4984_ (.D(_0331_),
    .CK(clknet_leaf_5_pclk),
    .Q(\mem[24] [9]),
    .QN(_2523_));
 DFF_X1 _4985_ (.D(_0332_),
    .CK(clknet_leaf_17_pclk),
    .Q(\mem[24] [10]),
    .QN(_2522_));
 DFF_X1 _4986_ (.D(_0333_),
    .CK(clknet_leaf_6_pclk),
    .Q(\mem[24] [11]),
    .QN(_2521_));
 DFF_X1 _4987_ (.D(_0334_),
    .CK(clknet_leaf_2_pclk),
    .Q(\mem[24] [12]),
    .QN(_2520_));
 DFF_X1 _4988_ (.D(_0335_),
    .CK(clknet_leaf_29_pclk),
    .Q(\mem[24] [13]),
    .QN(_2519_));
 DFF_X1 _4989_ (.D(_0336_),
    .CK(clknet_leaf_26_pclk),
    .Q(\mem[24] [14]),
    .QN(_2518_));
 DFF_X1 _4990_ (.D(_0337_),
    .CK(clknet_leaf_26_pclk),
    .Q(\mem[24] [15]),
    .QN(_2517_));
 DFF_X1 _4991_ (.D(_0338_),
    .CK(clknet_leaf_11_pclk),
    .Q(\mem[24] [16]),
    .QN(_2516_));
 DFF_X1 _4992_ (.D(_0339_),
    .CK(clknet_leaf_14_pclk),
    .Q(\mem[24] [17]),
    .QN(_2515_));
 DFF_X1 _4993_ (.D(_0340_),
    .CK(clknet_leaf_9_pclk),
    .Q(\mem[24] [18]),
    .QN(_2514_));
 DFF_X1 _4994_ (.D(_0341_),
    .CK(clknet_leaf_5_pclk),
    .Q(\mem[24] [19]),
    .QN(_2513_));
 DFF_X1 _4995_ (.D(_0342_),
    .CK(clknet_leaf_34_pclk),
    .Q(\mem[24] [20]),
    .QN(_2512_));
 DFF_X1 _4996_ (.D(_0343_),
    .CK(clknet_leaf_15_pclk),
    .Q(\mem[24] [21]),
    .QN(_2511_));
 DFF_X1 _4997_ (.D(_0344_),
    .CK(clknet_leaf_7_pclk),
    .Q(\mem[24] [22]),
    .QN(_2510_));
 DFF_X1 _4998_ (.D(_0345_),
    .CK(clknet_leaf_21_pclk),
    .Q(\mem[24] [23]),
    .QN(_2509_));
 DFF_X1 _4999_ (.D(_0346_),
    .CK(clknet_leaf_16_pclk),
    .Q(\mem[24] [24]),
    .QN(_2508_));
 DFF_X1 _5000_ (.D(_0347_),
    .CK(clknet_leaf_20_pclk),
    .Q(\mem[24] [25]),
    .QN(_2507_));
 DFF_X1 _5001_ (.D(_0348_),
    .CK(clknet_leaf_8_pclk),
    .Q(\mem[24] [26]),
    .QN(_2506_));
 DFF_X1 _5002_ (.D(_0349_),
    .CK(clknet_leaf_0_pclk),
    .Q(\mem[24] [27]),
    .QN(_2505_));
 DFF_X1 _5003_ (.D(_0350_),
    .CK(clknet_leaf_29_pclk),
    .Q(\mem[24] [28]),
    .QN(_2504_));
 DFF_X1 _5004_ (.D(_0351_),
    .CK(clknet_leaf_31_pclk),
    .Q(\mem[24] [29]),
    .QN(_2503_));
 DFF_X1 _5005_ (.D(_0352_),
    .CK(clknet_leaf_19_pclk),
    .Q(\mem[24] [30]),
    .QN(_2502_));
 DFF_X1 _5006_ (.D(_0353_),
    .CK(clknet_leaf_28_pclk),
    .Q(\mem[24] [31]),
    .QN(_2501_));
 DFF_X1 _5007_ (.D(_0354_),
    .CK(clknet_leaf_19_pclk),
    .Q(\mem[9] [0]),
    .QN(_2500_));
 DFF_X1 _5008_ (.D(_0355_),
    .CK(clknet_leaf_26_pclk),
    .Q(\mem[9] [1]),
    .QN(_2499_));
 DFF_X1 _5009_ (.D(_0356_),
    .CK(clknet_leaf_3_pclk),
    .Q(\mem[9] [2]),
    .QN(_2498_));
 DFF_X1 _5010_ (.D(_0357_),
    .CK(clknet_leaf_14_pclk),
    .Q(\mem[9] [3]),
    .QN(_2497_));
 DFF_X1 _5011_ (.D(_0358_),
    .CK(clknet_leaf_22_pclk),
    .Q(\mem[9] [4]),
    .QN(_2496_));
 DFF_X1 _5012_ (.D(_0359_),
    .CK(clknet_leaf_10_pclk),
    .Q(\mem[9] [5]),
    .QN(_2495_));
 DFF_X1 _5013_ (.D(_0360_),
    .CK(clknet_leaf_1_pclk),
    .Q(\mem[9] [6]),
    .QN(_2494_));
 DFF_X1 _5014_ (.D(_0361_),
    .CK(clknet_leaf_27_pclk),
    .Q(\mem[9] [7]),
    .QN(_2493_));
 DFF_X1 _5015_ (.D(_0362_),
    .CK(clknet_leaf_34_pclk),
    .Q(\mem[9] [8]),
    .QN(_2492_));
 DFF_X1 _5016_ (.D(_0363_),
    .CK(clknet_leaf_1_pclk),
    .Q(\mem[9] [9]),
    .QN(_2491_));
 DFF_X1 _5017_ (.D(_0364_),
    .CK(clknet_leaf_16_pclk),
    .Q(\mem[9] [10]),
    .QN(_2490_));
 DFF_X1 _5018_ (.D(_0365_),
    .CK(clknet_leaf_6_pclk),
    .Q(\mem[9] [11]),
    .QN(_2489_));
 DFF_X1 _5019_ (.D(_0366_),
    .CK(clknet_leaf_30_pclk),
    .Q(\mem[9] [12]),
    .QN(_2488_));
 DFF_X1 _5020_ (.D(_0367_),
    .CK(clknet_leaf_21_pclk),
    .Q(\mem[9] [13]),
    .QN(_2487_));
 DFF_X1 _5021_ (.D(_0368_),
    .CK(clknet_leaf_25_pclk),
    .Q(\mem[9] [14]),
    .QN(_2486_));
 DFF_X1 _5022_ (.D(_0369_),
    .CK(clknet_leaf_25_pclk),
    .Q(\mem[9] [15]),
    .QN(_2485_));
 DFF_X1 _5023_ (.D(_0370_),
    .CK(clknet_leaf_11_pclk),
    .Q(\mem[9] [16]),
    .QN(_2484_));
 DFF_X1 _5024_ (.D(_0371_),
    .CK(clknet_leaf_13_pclk),
    .Q(\mem[9] [17]),
    .QN(_2483_));
 DFF_X1 _5025_ (.D(_0372_),
    .CK(clknet_leaf_11_pclk),
    .Q(\mem[9] [18]),
    .QN(_2482_));
 DFF_X1 _5026_ (.D(_0373_),
    .CK(clknet_leaf_6_pclk),
    .Q(\mem[9] [19]),
    .QN(_2481_));
 DFF_X1 _5027_ (.D(_0374_),
    .CK(clknet_leaf_33_pclk),
    .Q(\mem[9] [20]),
    .QN(_2480_));
 DFF_X1 _5028_ (.D(_0375_),
    .CK(clknet_leaf_15_pclk),
    .Q(\mem[9] [21]),
    .QN(_2479_));
 DFF_X1 _5029_ (.D(_0376_),
    .CK(clknet_leaf_8_pclk),
    .Q(\mem[9] [22]),
    .QN(_2478_));
 DFF_X1 _5030_ (.D(_0377_),
    .CK(clknet_leaf_29_pclk),
    .Q(\mem[9] [23]),
    .QN(_2477_));
 DFF_X1 _5031_ (.D(_0378_),
    .CK(clknet_leaf_16_pclk),
    .Q(\mem[9] [24]),
    .QN(_2476_));
 DFF_X1 _5032_ (.D(_0379_),
    .CK(clknet_leaf_21_pclk),
    .Q(\mem[9] [25]),
    .QN(_2475_));
 DFF_X1 _5033_ (.D(_0380_),
    .CK(clknet_leaf_8_pclk),
    .Q(\mem[9] [26]),
    .QN(_2474_));
 DFF_X1 _5034_ (.D(_0381_),
    .CK(clknet_leaf_0_pclk),
    .Q(\mem[9] [27]),
    .QN(_2473_));
 DFF_X1 _5035_ (.D(_0382_),
    .CK(clknet_leaf_23_pclk),
    .Q(\mem[9] [28]),
    .QN(_2472_));
 DFF_X1 _5036_ (.D(_0383_),
    .CK(clknet_leaf_32_pclk),
    .Q(\mem[9] [29]),
    .QN(_2471_));
 DFF_X1 _5037_ (.D(_0384_),
    .CK(clknet_leaf_19_pclk),
    .Q(\mem[9] [30]),
    .QN(_2470_));
 DFF_X1 _5038_ (.D(_0385_),
    .CK(clknet_leaf_31_pclk),
    .Q(\mem[9] [31]),
    .QN(_2469_));
 DFF_X1 _5039_ (.D(_0386_),
    .CK(clknet_leaf_18_pclk),
    .Q(\mem[20] [0]),
    .QN(_2468_));
 DFF_X1 _5040_ (.D(_0387_),
    .CK(clknet_leaf_27_pclk),
    .Q(\mem[20] [1]),
    .QN(_2467_));
 DFF_X1 _5041_ (.D(_0388_),
    .CK(clknet_leaf_3_pclk),
    .Q(\mem[20] [2]),
    .QN(_2466_));
 DFF_X1 _5042_ (.D(_0389_),
    .CK(clknet_leaf_14_pclk),
    .Q(\mem[20] [3]),
    .QN(_2465_));
 DFF_X1 _5043_ (.D(_0390_),
    .CK(clknet_leaf_23_pclk),
    .Q(\mem[20] [4]),
    .QN(_2464_));
 DFF_X1 _5044_ (.D(_0391_),
    .CK(clknet_leaf_14_pclk),
    .Q(\mem[20] [5]),
    .QN(_2463_));
 DFF_X1 _5045_ (.D(_0392_),
    .CK(clknet_leaf_2_pclk),
    .Q(\mem[20] [6]),
    .QN(_2462_));
 DFF_X1 _5046_ (.D(_0393_),
    .CK(clknet_leaf_27_pclk),
    .Q(\mem[20] [7]),
    .QN(_2461_));
 DFF_X1 _5047_ (.D(_0394_),
    .CK(clknet_leaf_34_pclk),
    .Q(\mem[20] [8]),
    .QN(_2460_));
 DFF_X1 _5048_ (.D(_0395_),
    .CK(clknet_leaf_2_pclk),
    .Q(\mem[20] [9]),
    .QN(_2459_));
 DFF_X1 _5049_ (.D(_0396_),
    .CK(clknet_leaf_18_pclk),
    .Q(\mem[20] [10]),
    .QN(_2458_));
 DFF_X1 _5050_ (.D(_0397_),
    .CK(clknet_leaf_4_pclk),
    .Q(\mem[20] [11]),
    .QN(_2457_));
 DFF_X1 _5051_ (.D(_0398_),
    .CK(clknet_leaf_31_pclk),
    .Q(\mem[20] [12]),
    .QN(_2456_));
 DFF_X1 _5052_ (.D(_0399_),
    .CK(clknet_leaf_29_pclk),
    .Q(\mem[20] [13]),
    .QN(_2455_));
 DFF_X1 _5053_ (.D(_0400_),
    .CK(clknet_leaf_25_pclk),
    .Q(\mem[20] [14]),
    .QN(_2454_));
 DFF_X1 _5054_ (.D(_0401_),
    .CK(clknet_leaf_24_pclk),
    .Q(\mem[20] [15]),
    .QN(_2453_));
 DFF_X1 _5055_ (.D(_0402_),
    .CK(clknet_leaf_11_pclk),
    .Q(\mem[20] [16]),
    .QN(_2452_));
 DFF_X1 _5056_ (.D(_0403_),
    .CK(clknet_leaf_13_pclk),
    .Q(\mem[20] [17]),
    .QN(_2451_));
 DFF_X1 _5057_ (.D(_0404_),
    .CK(clknet_leaf_11_pclk),
    .Q(\mem[20] [18]),
    .QN(_2450_));
 DFF_X1 _5058_ (.D(_0405_),
    .CK(clknet_leaf_6_pclk),
    .Q(\mem[20] [19]),
    .QN(_2449_));
 DFF_X1 _5059_ (.D(_0406_),
    .CK(clknet_leaf_33_pclk),
    .Q(\mem[20] [20]),
    .QN(_2448_));
 DFF_X1 _5060_ (.D(_0407_),
    .CK(clknet_leaf_13_pclk),
    .Q(\mem[20] [21]),
    .QN(_2447_));
 DFF_X1 _5061_ (.D(_0408_),
    .CK(clknet_leaf_7_pclk),
    .Q(\mem[20] [22]),
    .QN(_2446_));
 DFF_X1 _5062_ (.D(_0409_),
    .CK(clknet_leaf_30_pclk),
    .Q(\mem[20] [23]),
    .QN(_2445_));
 DFF_X1 _5063_ (.D(_0410_),
    .CK(clknet_leaf_17_pclk),
    .Q(\mem[20] [24]),
    .QN(_2444_));
 DFF_X1 _5064_ (.D(_0411_),
    .CK(clknet_leaf_20_pclk),
    .Q(\mem[20] [25]),
    .QN(_2443_));
 DFF_X1 _5065_ (.D(_0412_),
    .CK(clknet_leaf_11_pclk),
    .Q(\mem[20] [26]),
    .QN(_2442_));
 DFF_X1 _5066_ (.D(_0413_),
    .CK(clknet_leaf_0_pclk),
    .Q(\mem[20] [27]),
    .QN(_2441_));
 DFF_X1 _5067_ (.D(_0414_),
    .CK(clknet_leaf_23_pclk),
    .Q(\mem[20] [28]),
    .QN(_2440_));
 DFF_X1 _5068_ (.D(_0415_),
    .CK(clknet_leaf_33_pclk),
    .Q(\mem[20] [29]),
    .QN(_2439_));
 DFF_X1 _5069_ (.D(_0416_),
    .CK(clknet_leaf_18_pclk),
    .Q(\mem[20] [30]),
    .QN(_2438_));
 DFF_X1 _5070_ (.D(_0417_),
    .CK(clknet_leaf_32_pclk),
    .Q(\mem[20] [31]),
    .QN(_2437_));
 DFF_X1 _5071_ (.D(_0418_),
    .CK(clknet_leaf_18_pclk),
    .Q(\mem[2] [0]),
    .QN(_2436_));
 DFF_X1 _5072_ (.D(_0419_),
    .CK(clknet_leaf_26_pclk),
    .Q(\mem[2] [1]),
    .QN(_2435_));
 DFF_X1 _5073_ (.D(_0420_),
    .CK(clknet_leaf_30_pclk),
    .Q(\mem[2] [2]),
    .QN(_2434_));
 DFF_X1 _5074_ (.D(_0421_),
    .CK(clknet_leaf_14_pclk),
    .Q(\mem[2] [3]),
    .QN(_2433_));
 DFF_X1 _5075_ (.D(_0422_),
    .CK(clknet_leaf_23_pclk),
    .Q(\mem[2] [4]),
    .QN(_2432_));
 DFF_X1 _5076_ (.D(_0423_),
    .CK(clknet_leaf_10_pclk),
    .Q(\mem[2] [5]),
    .QN(_2431_));
 DFF_X1 _5077_ (.D(_0424_),
    .CK(clknet_leaf_2_pclk),
    .Q(\mem[2] [6]),
    .QN(_2430_));
 DFF_X1 _5078_ (.D(_0425_),
    .CK(clknet_leaf_28_pclk),
    .Q(\mem[2] [7]),
    .QN(_2429_));
 DFF_X1 _5079_ (.D(_0426_),
    .CK(clknet_leaf_33_pclk),
    .Q(\mem[2] [8]),
    .QN(_2428_));
 DFF_X1 _5080_ (.D(_0427_),
    .CK(clknet_leaf_5_pclk),
    .Q(\mem[2] [9]),
    .QN(_2427_));
 DFF_X1 _5081_ (.D(_0428_),
    .CK(clknet_leaf_17_pclk),
    .Q(\mem[2] [10]),
    .QN(_2426_));
 DFF_X1 _5082_ (.D(_0429_),
    .CK(clknet_leaf_4_pclk),
    .Q(\mem[2] [11]),
    .QN(_2425_));
 DFF_X1 _5083_ (.D(_0430_),
    .CK(clknet_leaf_31_pclk),
    .Q(\mem[2] [12]),
    .QN(_2424_));
 DFF_X1 _5084_ (.D(_0431_),
    .CK(clknet_leaf_21_pclk),
    .Q(\mem[2] [13]),
    .QN(_2423_));
 DFF_X1 _5085_ (.D(_0432_),
    .CK(clknet_leaf_25_pclk),
    .Q(\mem[2] [14]),
    .QN(_2422_));
 DFF_X1 _5086_ (.D(_0433_),
    .CK(clknet_leaf_25_pclk),
    .Q(\mem[2] [15]),
    .QN(_2421_));
 DFF_X1 _5087_ (.D(_0434_),
    .CK(clknet_leaf_12_pclk),
    .Q(\mem[2] [16]),
    .QN(_2420_));
 DFF_X1 _5088_ (.D(_0435_),
    .CK(clknet_leaf_13_pclk),
    .Q(\mem[2] [17]),
    .QN(_2419_));
 DFF_X1 _5089_ (.D(_0436_),
    .CK(clknet_leaf_11_pclk),
    .Q(\mem[2] [18]),
    .QN(_2418_));
 DFF_X1 _5090_ (.D(_0437_),
    .CK(clknet_leaf_5_pclk),
    .Q(\mem[2] [19]),
    .QN(_2417_));
 DFF_X1 _5091_ (.D(_0438_),
    .CK(clknet_leaf_0_pclk),
    .Q(\mem[2] [20]),
    .QN(_2416_));
 DFF_X1 _5092_ (.D(_0439_),
    .CK(clknet_leaf_16_pclk),
    .Q(\mem[2] [21]),
    .QN(_2415_));
 DFF_X1 _5093_ (.D(_0440_),
    .CK(clknet_leaf_7_pclk),
    .Q(\mem[2] [22]),
    .QN(_2414_));
 DFF_X1 _5094_ (.D(_0441_),
    .CK(clknet_leaf_29_pclk),
    .Q(\mem[2] [23]),
    .QN(_2413_));
 DFF_X1 _5095_ (.D(_0442_),
    .CK(clknet_leaf_16_pclk),
    .Q(\mem[2] [24]),
    .QN(_2412_));
 DFF_X1 _5096_ (.D(_0443_),
    .CK(clknet_leaf_13_pclk),
    .Q(\mem[2] [25]),
    .QN(_2411_));
 DFF_X1 _5097_ (.D(_0444_),
    .CK(clknet_leaf_9_pclk),
    .Q(\mem[2] [26]),
    .QN(_2410_));
 DFF_X1 _5098_ (.D(_0445_),
    .CK(clknet_leaf_0_pclk),
    .Q(\mem[2] [27]),
    .QN(_2409_));
 DFF_X1 _5099_ (.D(_0446_),
    .CK(clknet_leaf_23_pclk),
    .Q(\mem[2] [28]),
    .QN(_2408_));
 DFF_X1 _5100_ (.D(_0447_),
    .CK(clknet_leaf_31_pclk),
    .Q(\mem[2] [29]),
    .QN(_2407_));
 DFF_X1 _5101_ (.D(_0448_),
    .CK(clknet_leaf_23_pclk),
    .Q(\mem[2] [30]),
    .QN(_2406_));
 DFF_X1 _5102_ (.D(_0449_),
    .CK(clknet_leaf_28_pclk),
    .Q(\mem[2] [31]),
    .QN(_2405_));
 DFF_X1 _5103_ (.D(_0450_),
    .CK(clknet_leaf_18_pclk),
    .Q(\mem[21] [0]),
    .QN(_2404_));
 DFF_X1 _5104_ (.D(_0451_),
    .CK(clknet_leaf_27_pclk),
    .Q(\mem[21] [1]),
    .QN(_2403_));
 DFF_X1 _5105_ (.D(_0452_),
    .CK(clknet_leaf_3_pclk),
    .Q(\mem[21] [2]),
    .QN(_2402_));
 DFF_X1 _5106_ (.D(_0453_),
    .CK(clknet_leaf_13_pclk),
    .Q(\mem[21] [3]),
    .QN(_2401_));
 DFF_X1 _5107_ (.D(_0454_),
    .CK(clknet_leaf_23_pclk),
    .Q(\mem[21] [4]),
    .QN(_2400_));
 DFF_X1 _5108_ (.D(_0455_),
    .CK(clknet_leaf_10_pclk),
    .Q(\mem[21] [5]),
    .QN(_2399_));
 DFF_X1 _5109_ (.D(_0456_),
    .CK(clknet_leaf_2_pclk),
    .Q(\mem[21] [6]),
    .QN(_2398_));
 DFF_X1 _5110_ (.D(_0457_),
    .CK(clknet_leaf_27_pclk),
    .Q(\mem[21] [7]),
    .QN(_2397_));
 DFF_X1 _5111_ (.D(_0458_),
    .CK(clknet_leaf_34_pclk),
    .Q(\mem[21] [8]),
    .QN(_2396_));
 DFF_X1 _5112_ (.D(_0459_),
    .CK(clknet_leaf_1_pclk),
    .Q(\mem[21] [9]),
    .QN(_2395_));
 DFF_X1 _5113_ (.D(_0460_),
    .CK(clknet_leaf_17_pclk),
    .Q(\mem[21] [10]),
    .QN(_2394_));
 DFF_X1 _5114_ (.D(_0461_),
    .CK(clknet_leaf_7_pclk),
    .Q(\mem[21] [11]),
    .QN(_2393_));
 DFF_X1 _5115_ (.D(_0462_),
    .CK(clknet_leaf_31_pclk),
    .Q(\mem[21] [12]),
    .QN(_2392_));
 DFF_X1 _5116_ (.D(_0463_),
    .CK(clknet_leaf_29_pclk),
    .Q(\mem[21] [13]),
    .QN(_2391_));
 DFF_X1 _5117_ (.D(_0464_),
    .CK(clknet_leaf_25_pclk),
    .Q(\mem[21] [14]),
    .QN(_2390_));
 DFF_X1 _5118_ (.D(_0465_),
    .CK(clknet_leaf_23_pclk),
    .Q(\mem[21] [15]),
    .QN(_2389_));
 DFF_X1 _5119_ (.D(_0466_),
    .CK(clknet_leaf_4_pclk),
    .Q(\mem[21] [16]),
    .QN(_2388_));
 DFF_X1 _5120_ (.D(_0467_),
    .CK(clknet_leaf_12_pclk),
    .Q(\mem[21] [17]),
    .QN(_2387_));
 DFF_X1 _5121_ (.D(_0468_),
    .CK(clknet_leaf_11_pclk),
    .Q(\mem[21] [18]),
    .QN(_2386_));
 DFF_X1 _5122_ (.D(_0469_),
    .CK(clknet_leaf_5_pclk),
    .Q(\mem[21] [19]),
    .QN(_2385_));
 DFF_X1 _5123_ (.D(_0470_),
    .CK(clknet_leaf_34_pclk),
    .Q(\mem[21] [20]),
    .QN(_2384_));
 DFF_X1 _5124_ (.D(_0471_),
    .CK(clknet_leaf_15_pclk),
    .Q(\mem[21] [21]),
    .QN(_2383_));
 DFF_X1 _5125_ (.D(_0472_),
    .CK(clknet_leaf_7_pclk),
    .Q(\mem[21] [22]),
    .QN(_2382_));
 DFF_X1 _5126_ (.D(_0473_),
    .CK(clknet_leaf_30_pclk),
    .Q(\mem[21] [23]),
    .QN(_2381_));
 DFF_X1 _5127_ (.D(_0474_),
    .CK(clknet_leaf_17_pclk),
    .Q(\mem[21] [24]),
    .QN(_2380_));
 DFF_X1 _5128_ (.D(_0475_),
    .CK(clknet_leaf_20_pclk),
    .Q(\mem[21] [25]),
    .QN(_2379_));
 DFF_X1 _5129_ (.D(_0476_),
    .CK(clknet_leaf_7_pclk),
    .Q(\mem[21] [26]),
    .QN(_2378_));
 DFF_X1 _5130_ (.D(_0477_),
    .CK(clknet_leaf_1_pclk),
    .Q(\mem[21] [27]),
    .QN(_2377_));
 DFF_X1 _5131_ (.D(_0478_),
    .CK(clknet_leaf_29_pclk),
    .Q(\mem[21] [28]),
    .QN(_2376_));
 DFF_X1 _5132_ (.D(_0479_),
    .CK(clknet_leaf_32_pclk),
    .Q(\mem[21] [29]),
    .QN(_2375_));
 DFF_X1 _5133_ (.D(_0480_),
    .CK(clknet_leaf_19_pclk),
    .Q(\mem[21] [30]),
    .QN(_2374_));
 DFF_X1 _5134_ (.D(_0481_),
    .CK(clknet_leaf_28_pclk),
    .Q(\mem[21] [31]),
    .QN(_2373_));
 DFF_X1 _5135_ (.D(_0482_),
    .CK(clknet_leaf_20_pclk),
    .Q(\mem[30] [0]),
    .QN(_2372_));
 DFF_X1 _5136_ (.D(_0483_),
    .CK(clknet_leaf_26_pclk),
    .Q(\mem[30] [1]),
    .QN(_2371_));
 DFF_X1 _5137_ (.D(_0484_),
    .CK(clknet_leaf_4_pclk),
    .Q(\mem[30] [2]),
    .QN(_2370_));
 DFF_X1 _5138_ (.D(_0485_),
    .CK(clknet_leaf_14_pclk),
    .Q(\mem[30] [3]),
    .QN(_2369_));
 DFF_X1 _5139_ (.D(_0486_),
    .CK(clknet_leaf_22_pclk),
    .Q(\mem[30] [4]),
    .QN(_2368_));
 DFF_X1 _5140_ (.D(_0487_),
    .CK(clknet_leaf_9_pclk),
    .Q(\mem[30] [5]),
    .QN(_2367_));
 DFF_X1 _5141_ (.D(_0488_),
    .CK(clknet_leaf_1_pclk),
    .Q(\mem[30] [6]),
    .QN(_2366_));
 DFF_X1 _5142_ (.D(_0489_),
    .CK(clknet_leaf_28_pclk),
    .Q(\mem[30] [7]),
    .QN(_2365_));
 DFF_X1 _5143_ (.D(_0490_),
    .CK(clknet_leaf_34_pclk),
    .Q(\mem[30] [8]),
    .QN(_2364_));
 DFF_X1 _5144_ (.D(_0491_),
    .CK(clknet_leaf_5_pclk),
    .Q(\mem[30] [9]),
    .QN(_2363_));
 DFF_X1 _5145_ (.D(_0492_),
    .CK(clknet_leaf_17_pclk),
    .Q(\mem[30] [10]),
    .QN(_2362_));
 DFF_X1 _5146_ (.D(_0493_),
    .CK(clknet_leaf_5_pclk),
    .Q(\mem[30] [11]),
    .QN(_2361_));
 DFF_X1 _5147_ (.D(_0494_),
    .CK(clknet_leaf_31_pclk),
    .Q(\mem[30] [12]),
    .QN(_2360_));
 DFF_X1 _5148_ (.D(_0495_),
    .CK(clknet_leaf_29_pclk),
    .Q(\mem[30] [13]),
    .QN(_2359_));
 DFF_X1 _5149_ (.D(_0496_),
    .CK(clknet_leaf_26_pclk),
    .Q(\mem[30] [14]),
    .QN(_2358_));
 DFF_X1 _5150_ (.D(_0497_),
    .CK(clknet_leaf_24_pclk),
    .Q(\mem[30] [15]),
    .QN(_2357_));
 DFF_X1 _5151_ (.D(_0498_),
    .CK(clknet_leaf_12_pclk),
    .Q(\mem[30] [16]),
    .QN(_2356_));
 DFF_X1 _5152_ (.D(_0499_),
    .CK(clknet_leaf_14_pclk),
    .Q(\mem[30] [17]),
    .QN(_2355_));
 DFF_X1 _5153_ (.D(_0500_),
    .CK(clknet_leaf_8_pclk),
    .Q(\mem[30] [18]),
    .QN(_2354_));
 DFF_X1 _5154_ (.D(_0501_),
    .CK(clknet_leaf_6_pclk),
    .Q(\mem[30] [19]),
    .QN(_2353_));
 DFF_X1 _5155_ (.D(_0502_),
    .CK(clknet_leaf_33_pclk),
    .Q(\mem[30] [20]),
    .QN(_2352_));
 DFF_X1 _5156_ (.D(_0503_),
    .CK(clknet_leaf_13_pclk),
    .Q(\mem[30] [21]),
    .QN(_2351_));
 DFF_X1 _5157_ (.D(_0504_),
    .CK(clknet_leaf_7_pclk),
    .Q(\mem[30] [22]),
    .QN(_2350_));
 DFF_X1 _5158_ (.D(_0505_),
    .CK(clknet_leaf_30_pclk),
    .Q(\mem[30] [23]),
    .QN(_2349_));
 DFF_X1 _5159_ (.D(_0506_),
    .CK(clknet_leaf_16_pclk),
    .Q(\mem[30] [24]),
    .QN(_2348_));
 DFF_X1 _5160_ (.D(_0507_),
    .CK(clknet_leaf_20_pclk),
    .Q(\mem[30] [25]),
    .QN(_2347_));
 DFF_X1 _5161_ (.D(_0508_),
    .CK(clknet_leaf_8_pclk),
    .Q(\mem[30] [26]),
    .QN(_2346_));
 DFF_X1 _5162_ (.D(_0509_),
    .CK(clknet_leaf_35_pclk),
    .Q(\mem[30] [27]),
    .QN(_2345_));
 DFF_X1 _5163_ (.D(_0510_),
    .CK(clknet_leaf_22_pclk),
    .Q(\mem[30] [28]),
    .QN(_2344_));
 DFF_X1 _5164_ (.D(_0511_),
    .CK(clknet_leaf_31_pclk),
    .Q(\mem[30] [29]),
    .QN(_2343_));
 DFF_X1 _5165_ (.D(_0512_),
    .CK(clknet_leaf_22_pclk),
    .Q(\mem[30] [30]),
    .QN(_2342_));
 DFF_X1 _5166_ (.D(_0513_),
    .CK(clknet_leaf_28_pclk),
    .Q(\mem[30] [31]),
    .QN(_2341_));
 DFF_X1 _5167_ (.D(_0514_),
    .CK(clknet_leaf_18_pclk),
    .Q(\mem[22] [0]),
    .QN(_2340_));
 DFF_X1 _5168_ (.D(_0515_),
    .CK(clknet_leaf_25_pclk),
    .Q(\mem[22] [1]),
    .QN(_2339_));
 DFF_X1 _5169_ (.D(_0516_),
    .CK(clknet_leaf_12_pclk),
    .Q(\mem[22] [2]),
    .QN(_2338_));
 DFF_X1 _5170_ (.D(_0517_),
    .CK(clknet_leaf_13_pclk),
    .Q(\mem[22] [3]),
    .QN(_2337_));
 DFF_X1 _5171_ (.D(_0518_),
    .CK(clknet_leaf_23_pclk),
    .Q(\mem[22] [4]),
    .QN(_2336_));
 DFF_X1 _5172_ (.D(_0519_),
    .CK(clknet_leaf_10_pclk),
    .Q(\mem[22] [5]),
    .QN(_2335_));
 DFF_X1 _5173_ (.D(_0520_),
    .CK(clknet_leaf_2_pclk),
    .Q(\mem[22] [6]),
    .QN(_2334_));
 DFF_X1 _5174_ (.D(_0521_),
    .CK(clknet_leaf_27_pclk),
    .Q(\mem[22] [7]),
    .QN(_2333_));
 DFF_X1 _5175_ (.D(_0522_),
    .CK(clknet_leaf_34_pclk),
    .Q(\mem[22] [8]),
    .QN(_2332_));
 DFF_X1 _5176_ (.D(_0523_),
    .CK(clknet_leaf_2_pclk),
    .Q(\mem[22] [9]),
    .QN(_2331_));
 DFF_X1 _5177_ (.D(_0524_),
    .CK(clknet_leaf_17_pclk),
    .Q(\mem[22] [10]),
    .QN(_2330_));
 DFF_X1 _5178_ (.D(_0525_),
    .CK(clknet_leaf_4_pclk),
    .Q(\mem[22] [11]),
    .QN(_2329_));
 DFF_X1 _5179_ (.D(_0526_),
    .CK(clknet_leaf_31_pclk),
    .Q(\mem[22] [12]),
    .QN(_2328_));
 DFF_X1 _5180_ (.D(_0527_),
    .CK(clknet_leaf_22_pclk),
    .Q(\mem[22] [13]),
    .QN(_2327_));
 DFF_X1 _5181_ (.D(_0528_),
    .CK(clknet_leaf_25_pclk),
    .Q(\mem[22] [14]),
    .QN(_2326_));
 DFF_X1 _5182_ (.D(_0529_),
    .CK(clknet_leaf_24_pclk),
    .Q(\mem[22] [15]),
    .QN(_2325_));
 DFF_X1 _5183_ (.D(_0530_),
    .CK(clknet_leaf_11_pclk),
    .Q(\mem[22] [16]),
    .QN(_2324_));
 DFF_X1 _5184_ (.D(_0531_),
    .CK(clknet_leaf_10_pclk),
    .Q(\mem[22] [17]),
    .QN(_2323_));
 DFF_X1 _5185_ (.D(_0532_),
    .CK(clknet_leaf_11_pclk),
    .Q(\mem[22] [18]),
    .QN(_2322_));
 DFF_X1 _5186_ (.D(_0533_),
    .CK(clknet_leaf_6_pclk),
    .Q(\mem[22] [19]),
    .QN(_2321_));
 DFF_X1 _5187_ (.D(_0534_),
    .CK(clknet_leaf_33_pclk),
    .Q(\mem[22] [20]),
    .QN(_2320_));
 DFF_X1 _5188_ (.D(_0535_),
    .CK(clknet_leaf_13_pclk),
    .Q(\mem[22] [21]),
    .QN(_2319_));
 DFF_X1 _5189_ (.D(_0536_),
    .CK(clknet_leaf_7_pclk),
    .Q(\mem[22] [22]),
    .QN(_2318_));
 DFF_X1 _5190_ (.D(_0537_),
    .CK(clknet_leaf_30_pclk),
    .Q(\mem[22] [23]),
    .QN(_2317_));
 DFF_X1 _5191_ (.D(_0538_),
    .CK(clknet_leaf_17_pclk),
    .Q(\mem[22] [24]),
    .QN(_2316_));
 DFF_X1 _5192_ (.D(_0539_),
    .CK(clknet_leaf_21_pclk),
    .Q(\mem[22] [25]),
    .QN(_2315_));
 DFF_X1 _5193_ (.D(_0540_),
    .CK(clknet_leaf_11_pclk),
    .Q(\mem[22] [26]),
    .QN(_2314_));
 DFF_X1 _5194_ (.D(_0541_),
    .CK(clknet_leaf_0_pclk),
    .Q(\mem[22] [27]),
    .QN(_2313_));
 DFF_X1 _5195_ (.D(_0542_),
    .CK(clknet_leaf_24_pclk),
    .Q(\mem[22] [28]),
    .QN(_2312_));
 DFF_X1 _5196_ (.D(_0543_),
    .CK(clknet_leaf_33_pclk),
    .Q(\mem[22] [29]),
    .QN(_2311_));
 DFF_X1 _5197_ (.D(_0544_),
    .CK(clknet_leaf_18_pclk),
    .Q(\mem[22] [30]),
    .QN(_2310_));
 DFF_X1 _5198_ (.D(_0545_),
    .CK(clknet_leaf_32_pclk),
    .Q(\mem[22] [31]),
    .QN(_2309_));
 DFFR_X1 _5199_ (.D(_0546_),
    .RN(prst_n),
    .CK(clknet_leaf_18_pclk),
    .Q(prdata[0]),
    .QN(_2308_));
 DFFR_X1 _5200_ (.D(_0547_),
    .RN(prst_n),
    .CK(clknet_leaf_25_pclk),
    .Q(prdata[1]),
    .QN(_2307_));
 DFFR_X2 _5201_ (.D(_0548_),
    .RN(prst_n),
    .CK(clknet_leaf_21_pclk),
    .Q(prdata[2]),
    .QN(_2306_));
 DFFR_X1 _5202_ (.D(_0549_),
    .RN(prst_n),
    .CK(clknet_leaf_14_pclk),
    .Q(prdata[3]),
    .QN(_2305_));
 DFFR_X1 _5203_ (.D(_0550_),
    .RN(prst_n),
    .CK(clknet_leaf_22_pclk),
    .Q(prdata[4]),
    .QN(_2304_));
 DFFR_X1 _5204_ (.D(_0551_),
    .RN(prst_n),
    .CK(clknet_leaf_10_pclk),
    .Q(prdata[5]),
    .QN(_2303_));
 DFFR_X1 _5205_ (.D(_0552_),
    .RN(prst_n),
    .CK(clknet_leaf_1_pclk),
    .Q(prdata[6]),
    .QN(_2302_));
 DFFR_X1 _5206_ (.D(_0553_),
    .RN(prst_n),
    .CK(clknet_leaf_28_pclk),
    .Q(prdata[7]),
    .QN(_2301_));
 DFFR_X1 _5207_ (.D(_0554_),
    .RN(prst_n),
    .CK(clknet_leaf_35_pclk),
    .Q(prdata[8]),
    .QN(_2300_));
 DFFR_X1 _5208_ (.D(_0555_),
    .RN(prst_n),
    .CK(clknet_leaf_1_pclk),
    .Q(prdata[9]),
    .QN(_2299_));
 DFFR_X1 _5209_ (.D(_0556_),
    .RN(prst_n),
    .CK(clknet_leaf_18_pclk),
    .Q(prdata[10]),
    .QN(_2298_));
 DFFR_X2 _5210_ (.D(_0557_),
    .RN(prst_n),
    .CK(clknet_leaf_6_pclk),
    .Q(prdata[11]),
    .QN(_2297_));
 DFFR_X2 _5211_ (.D(_0558_),
    .RN(prst_n),
    .CK(clknet_leaf_30_pclk),
    .Q(prdata[12]),
    .QN(_2296_));
 DFFR_X2 _5212_ (.D(_0559_),
    .RN(prst_n),
    .CK(clknet_leaf_22_pclk),
    .Q(prdata[13]),
    .QN(_2295_));
 DFFR_X1 _5213_ (.D(_0560_),
    .RN(prst_n),
    .CK(clknet_leaf_25_pclk),
    .Q(prdata[14]),
    .QN(_2294_));
 DFFR_X1 _5214_ (.D(_0561_),
    .RN(prst_n),
    .CK(clknet_leaf_24_pclk),
    .Q(prdata[15]),
    .QN(_2293_));
 DFFR_X2 _5215_ (.D(_0562_),
    .RN(prst_n),
    .CK(clknet_leaf_3_pclk),
    .Q(prdata[16]),
    .QN(_2292_));
 DFFR_X2 _5216_ (.D(_0563_),
    .RN(prst_n),
    .CK(clknet_leaf_12_pclk),
    .Q(prdata[17]),
    .QN(_2291_));
 DFFR_X1 _5217_ (.D(_0564_),
    .RN(prst_n),
    .CK(clknet_leaf_9_pclk),
    .Q(prdata[18]),
    .QN(_2290_));
 DFFR_X1 _5218_ (.D(_0565_),
    .RN(prst_n),
    .CK(clknet_leaf_5_pclk),
    .Q(prdata[19]),
    .QN(_2289_));
 DFFR_X1 _5219_ (.D(_0566_),
    .RN(prst_n),
    .CK(clknet_leaf_34_pclk),
    .Q(prdata[20]),
    .QN(_2288_));
 DFFR_X1 _5220_ (.D(_0567_),
    .RN(prst_n),
    .CK(clknet_leaf_15_pclk),
    .Q(prdata[21]),
    .QN(_2287_));
 DFFR_X1 _5221_ (.D(_0568_),
    .RN(prst_n),
    .CK(clknet_leaf_7_pclk),
    .Q(prdata[22]),
    .QN(_2286_));
 DFFR_X2 _5222_ (.D(_0569_),
    .RN(prst_n),
    .CK(clknet_leaf_21_pclk),
    .Q(prdata[23]),
    .QN(_2285_));
 DFFR_X1 _5223_ (.D(_0570_),
    .RN(prst_n),
    .CK(clknet_leaf_17_pclk),
    .Q(prdata[24]),
    .QN(_2284_));
 DFFR_X1 _5224_ (.D(_0571_),
    .RN(prst_n),
    .CK(clknet_leaf_5_pclk),
    .Q(prdata[25]),
    .QN(_2283_));
 DFFR_X1 _5225_ (.D(_0572_),
    .RN(prst_n),
    .CK(clknet_leaf_8_pclk),
    .Q(prdata[26]),
    .QN(_2282_));
 DFFR_X1 _5226_ (.D(_0573_),
    .RN(prst_n),
    .CK(clknet_leaf_0_pclk),
    .Q(prdata[27]),
    .QN(_2281_));
 DFFR_X1 _5227_ (.D(_0574_),
    .RN(prst_n),
    .CK(clknet_leaf_23_pclk),
    .Q(prdata[28]),
    .QN(_2280_));
 DFFR_X1 _5228_ (.D(_0575_),
    .RN(prst_n),
    .CK(clknet_leaf_32_pclk),
    .Q(prdata[29]),
    .QN(_2279_));
 DFFR_X1 _5229_ (.D(_0576_),
    .RN(prst_n),
    .CK(clknet_leaf_19_pclk),
    .Q(prdata[30]),
    .QN(_2278_));
 DFFR_X2 _5230_ (.D(_0577_),
    .RN(prst_n),
    .CK(clknet_leaf_28_pclk),
    .Q(prdata[31]),
    .QN(_2277_));
 DFF_X1 _5231_ (.D(_0578_),
    .CK(clknet_leaf_20_pclk),
    .Q(\mem[1] [0]),
    .QN(_2276_));
 DFF_X1 _5232_ (.D(_0579_),
    .CK(clknet_leaf_26_pclk),
    .Q(\mem[1] [1]),
    .QN(_2275_));
 DFF_X1 _5233_ (.D(_0580_),
    .CK(clknet_leaf_3_pclk),
    .Q(\mem[1] [2]),
    .QN(_2274_));
 DFF_X1 _5234_ (.D(_0581_),
    .CK(clknet_leaf_14_pclk),
    .Q(\mem[1] [3]),
    .QN(_2273_));
 DFF_X1 _5235_ (.D(_0582_),
    .CK(clknet_leaf_23_pclk),
    .Q(\mem[1] [4]),
    .QN(_2272_));
 DFF_X1 _5236_ (.D(_0583_),
    .CK(clknet_leaf_14_pclk),
    .Q(\mem[1] [5]),
    .QN(_2271_));
 DFF_X1 _5237_ (.D(_0584_),
    .CK(clknet_leaf_0_pclk),
    .Q(\mem[1] [6]),
    .QN(_2270_));
 DFF_X1 _5238_ (.D(_0585_),
    .CK(clknet_leaf_28_pclk),
    .Q(\mem[1] [7]),
    .QN(_2269_));
 DFF_X1 _5239_ (.D(_0586_),
    .CK(clknet_leaf_0_pclk),
    .Q(\mem[1] [8]),
    .QN(_2268_));
 DFF_X1 _5240_ (.D(_0587_),
    .CK(clknet_leaf_4_pclk),
    .Q(\mem[1] [9]),
    .QN(_2267_));
 DFF_X1 _5241_ (.D(_0588_),
    .CK(clknet_leaf_17_pclk),
    .Q(\mem[1] [10]),
    .QN(_2266_));
 DFF_X1 _5242_ (.D(_0589_),
    .CK(clknet_leaf_6_pclk),
    .Q(\mem[1] [11]),
    .QN(_2265_));
 DFF_X1 _5243_ (.D(_0590_),
    .CK(clknet_leaf_2_pclk),
    .Q(\mem[1] [12]),
    .QN(_2264_));
 DFF_X1 _5244_ (.D(_0591_),
    .CK(clknet_leaf_21_pclk),
    .Q(\mem[1] [13]),
    .QN(_2263_));
 DFF_X1 _5245_ (.D(_0592_),
    .CK(clknet_leaf_25_pclk),
    .Q(\mem[1] [14]),
    .QN(_2262_));
 DFF_X1 _5246_ (.D(_0593_),
    .CK(clknet_leaf_25_pclk),
    .Q(\mem[1] [15]),
    .QN(_2261_));
 DFF_X1 _5247_ (.D(_0594_),
    .CK(clknet_leaf_12_pclk),
    .Q(\mem[1] [16]),
    .QN(_2260_));
 DFF_X1 _5248_ (.D(_0595_),
    .CK(clknet_leaf_12_pclk),
    .Q(\mem[1] [17]),
    .QN(_2259_));
 DFF_X1 _5249_ (.D(_0596_),
    .CK(clknet_leaf_11_pclk),
    .Q(\mem[1] [18]),
    .QN(_2258_));
 DFF_X1 _5250_ (.D(_0597_),
    .CK(clknet_leaf_4_pclk),
    .Q(\mem[1] [19]),
    .QN(_2257_));
 DFF_X1 _5251_ (.D(_0598_),
    .CK(clknet_leaf_33_pclk),
    .Q(\mem[1] [20]),
    .QN(_2256_));
 DFF_X1 _5252_ (.D(_0599_),
    .CK(clknet_leaf_16_pclk),
    .Q(\mem[1] [21]),
    .QN(_2255_));
 DFF_X1 _5253_ (.D(_0600_),
    .CK(clknet_leaf_9_pclk),
    .Q(\mem[1] [22]),
    .QN(_2254_));
 DFF_X1 _5254_ (.D(_0601_),
    .CK(clknet_leaf_30_pclk),
    .Q(\mem[1] [23]),
    .QN(_2253_));
 DFF_X1 _5255_ (.D(_0602_),
    .CK(clknet_leaf_16_pclk),
    .Q(\mem[1] [24]),
    .QN(_2252_));
 DFF_X1 _5256_ (.D(_0603_),
    .CK(clknet_leaf_12_pclk),
    .Q(\mem[1] [25]),
    .QN(_2251_));
 DFF_X1 _5257_ (.D(_0604_),
    .CK(clknet_leaf_9_pclk),
    .Q(\mem[1] [26]),
    .QN(_2250_));
 DFF_X1 _5258_ (.D(_0605_),
    .CK(clknet_leaf_0_pclk),
    .Q(\mem[1] [27]),
    .QN(_2249_));
 DFF_X1 _5259_ (.D(_0606_),
    .CK(clknet_leaf_23_pclk),
    .Q(\mem[1] [28]),
    .QN(_2248_));
 DFF_X1 _5260_ (.D(_0607_),
    .CK(clknet_leaf_32_pclk),
    .Q(\mem[1] [29]),
    .QN(_2247_));
 DFF_X1 _5261_ (.D(_0608_),
    .CK(clknet_leaf_19_pclk),
    .Q(\mem[1] [30]),
    .QN(_2246_));
 DFF_X1 _5262_ (.D(_0609_),
    .CK(clknet_leaf_28_pclk),
    .Q(\mem[1] [31]),
    .QN(_2245_));
 DFF_X1 _5263_ (.D(_0610_),
    .CK(clknet_leaf_18_pclk),
    .Q(\mem[23] [0]),
    .QN(_2244_));
 DFF_X1 _5264_ (.D(_0611_),
    .CK(clknet_leaf_26_pclk),
    .Q(\mem[23] [1]),
    .QN(_2243_));
 DFF_X1 _5265_ (.D(_0612_),
    .CK(clknet_leaf_12_pclk),
    .Q(\mem[23] [2]),
    .QN(_2242_));
 DFF_X1 _5266_ (.D(_0613_),
    .CK(clknet_leaf_14_pclk),
    .Q(\mem[23] [3]),
    .QN(_2241_));
 DFF_X1 _5267_ (.D(_0614_),
    .CK(clknet_leaf_23_pclk),
    .Q(\mem[23] [4]),
    .QN(_2240_));
 DFF_X1 _5268_ (.D(_0615_),
    .CK(clknet_leaf_10_pclk),
    .Q(\mem[23] [5]),
    .QN(_2239_));
 DFF_X1 _5269_ (.D(_0616_),
    .CK(clknet_leaf_1_pclk),
    .Q(\mem[23] [6]),
    .QN(_2238_));
 DFF_X1 _5270_ (.D(_0617_),
    .CK(clknet_leaf_28_pclk),
    .Q(\mem[23] [7]),
    .QN(_2237_));
 DFF_X1 _5271_ (.D(_0618_),
    .CK(clknet_leaf_34_pclk),
    .Q(\mem[23] [8]),
    .QN(_2236_));
 DFF_X1 _5272_ (.D(_0619_),
    .CK(clknet_leaf_1_pclk),
    .Q(\mem[23] [9]),
    .QN(_2235_));
 DFF_X1 _5273_ (.D(_0620_),
    .CK(clknet_leaf_18_pclk),
    .Q(\mem[23] [10]),
    .QN(_2234_));
 DFF_X1 _5274_ (.D(_0621_),
    .CK(clknet_leaf_4_pclk),
    .Q(\mem[23] [11]),
    .QN(_2233_));
 DFF_X1 _5275_ (.D(_0622_),
    .CK(clknet_leaf_30_pclk),
    .Q(\mem[23] [12]),
    .QN(_2232_));
 DFF_X1 _5276_ (.D(_0623_),
    .CK(clknet_leaf_22_pclk),
    .Q(\mem[23] [13]),
    .QN(_2231_));
 DFF_X1 _5277_ (.D(_0624_),
    .CK(clknet_leaf_25_pclk),
    .Q(\mem[23] [14]),
    .QN(_2230_));
 DFF_X1 _5278_ (.D(_0625_),
    .CK(clknet_leaf_24_pclk),
    .Q(\mem[23] [15]),
    .QN(_2229_));
 DFF_X1 _5279_ (.D(_0626_),
    .CK(clknet_leaf_11_pclk),
    .Q(\mem[23] [16]),
    .QN(_2228_));
 DFF_X1 _5280_ (.D(_0627_),
    .CK(clknet_leaf_11_pclk),
    .Q(\mem[23] [17]),
    .QN(_2227_));
 DFF_X1 _5281_ (.D(_0628_),
    .CK(clknet_leaf_9_pclk),
    .Q(\mem[23] [18]),
    .QN(_2226_));
 DFF_X1 _5282_ (.D(_0629_),
    .CK(clknet_leaf_5_pclk),
    .Q(\mem[23] [19]),
    .QN(_2225_));
 DFF_X1 _5283_ (.D(_0630_),
    .CK(clknet_leaf_34_pclk),
    .Q(\mem[23] [20]),
    .QN(_2224_));
 DFF_X1 _5284_ (.D(_0631_),
    .CK(clknet_leaf_13_pclk),
    .Q(\mem[23] [21]),
    .QN(_2223_));
 DFF_X1 _5285_ (.D(_0632_),
    .CK(clknet_leaf_7_pclk),
    .Q(\mem[23] [22]),
    .QN(_2222_));
 DFF_X1 _5286_ (.D(_0633_),
    .CK(clknet_leaf_30_pclk),
    .Q(\mem[23] [23]),
    .QN(_2221_));
 DFF_X1 _5287_ (.D(_0634_),
    .CK(clknet_leaf_17_pclk),
    .Q(\mem[23] [24]),
    .QN(_2220_));
 DFF_X1 _5288_ (.D(_0635_),
    .CK(clknet_leaf_12_pclk),
    .Q(\mem[23] [25]),
    .QN(_2219_));
 DFF_X1 _5289_ (.D(_0636_),
    .CK(clknet_leaf_7_pclk),
    .Q(\mem[23] [26]),
    .QN(_2218_));
 DFF_X1 _5290_ (.D(_0637_),
    .CK(clknet_leaf_1_pclk),
    .Q(\mem[23] [27]),
    .QN(_2217_));
 DFF_X1 _5291_ (.D(_0638_),
    .CK(clknet_leaf_22_pclk),
    .Q(\mem[23] [28]),
    .QN(_2216_));
 DFF_X1 _5292_ (.D(_0639_),
    .CK(clknet_leaf_32_pclk),
    .Q(\mem[23] [29]),
    .QN(_2215_));
 DFF_X1 _5293_ (.D(_0640_),
    .CK(clknet_leaf_19_pclk),
    .Q(\mem[23] [30]),
    .QN(_2214_));
 DFF_X1 _5294_ (.D(_0641_),
    .CK(clknet_leaf_28_pclk),
    .Q(\mem[23] [31]),
    .QN(_2213_));
 DFF_X1 _5295_ (.D(_0642_),
    .CK(clknet_leaf_18_pclk),
    .Q(\mem[25] [0]),
    .QN(_2212_));
 DFF_X1 _5296_ (.D(_0643_),
    .CK(clknet_leaf_27_pclk),
    .Q(\mem[25] [1]),
    .QN(_2211_));
 DFF_X1 _5297_ (.D(_0644_),
    .CK(clknet_leaf_3_pclk),
    .Q(\mem[25] [2]),
    .QN(_2210_));
 DFF_X1 _5298_ (.D(_0645_),
    .CK(clknet_leaf_14_pclk),
    .Q(\mem[25] [3]),
    .QN(_2209_));
 DFF_X1 _5299_ (.D(_0646_),
    .CK(clknet_leaf_22_pclk),
    .Q(\mem[25] [4]),
    .QN(_2208_));
 DFF_X1 _5300_ (.D(_0647_),
    .CK(clknet_leaf_10_pclk),
    .Q(\mem[25] [5]),
    .QN(_2207_));
 DFF_X1 _5301_ (.D(_0648_),
    .CK(clknet_leaf_0_pclk),
    .Q(\mem[25] [6]),
    .QN(_2206_));
 DFF_X1 _5302_ (.D(_0649_),
    .CK(clknet_leaf_28_pclk),
    .Q(\mem[25] [7]),
    .QN(_2205_));
 DFF_X1 _5303_ (.D(_0650_),
    .CK(clknet_leaf_34_pclk),
    .Q(\mem[25] [8]),
    .QN(_2204_));
 DFF_X1 _5304_ (.D(_0651_),
    .CK(clknet_leaf_1_pclk),
    .Q(\mem[25] [9]),
    .QN(_2203_));
 DFF_X1 _5305_ (.D(_0652_),
    .CK(clknet_leaf_17_pclk),
    .Q(\mem[25] [10]),
    .QN(_2202_));
 DFF_X1 _5306_ (.D(_0653_),
    .CK(clknet_leaf_7_pclk),
    .Q(\mem[25] [11]),
    .QN(_2201_));
 DFF_X1 _5307_ (.D(_0654_),
    .CK(clknet_leaf_2_pclk),
    .Q(\mem[25] [12]),
    .QN(_2200_));
 DFF_X1 _5308_ (.D(_0655_),
    .CK(clknet_leaf_22_pclk),
    .Q(\mem[25] [13]),
    .QN(_2199_));
 DFF_X1 _5309_ (.D(_0656_),
    .CK(clknet_leaf_25_pclk),
    .Q(\mem[25] [14]),
    .QN(_2198_));
 DFF_X1 _5310_ (.D(_0657_),
    .CK(clknet_leaf_24_pclk),
    .Q(\mem[25] [15]),
    .QN(_2197_));
 DFF_X1 _5311_ (.D(_0658_),
    .CK(clknet_leaf_11_pclk),
    .Q(\mem[25] [16]),
    .QN(_2196_));
 DFF_X1 _5312_ (.D(_0659_),
    .CK(clknet_leaf_13_pclk),
    .Q(\mem[25] [17]),
    .QN(_2195_));
 DFF_X1 _5313_ (.D(_0660_),
    .CK(clknet_leaf_11_pclk),
    .Q(\mem[25] [18]),
    .QN(_2194_));
 DFF_X1 _5314_ (.D(_0661_),
    .CK(clknet_leaf_6_pclk),
    .Q(\mem[25] [19]),
    .QN(_2193_));
 DFF_X1 _5315_ (.D(_0662_),
    .CK(clknet_leaf_34_pclk),
    .Q(\mem[25] [20]),
    .QN(_2192_));
 DFF_X1 _5316_ (.D(_0663_),
    .CK(clknet_leaf_15_pclk),
    .Q(\mem[25] [21]),
    .QN(_2191_));
 DFF_X1 _5317_ (.D(_0664_),
    .CK(clknet_leaf_7_pclk),
    .Q(\mem[25] [22]),
    .QN(_2190_));
 DFF_X1 _5318_ (.D(_0665_),
    .CK(clknet_leaf_21_pclk),
    .Q(\mem[25] [23]),
    .QN(_2189_));
 DFF_X1 _5319_ (.D(_0666_),
    .CK(clknet_leaf_16_pclk),
    .Q(\mem[25] [24]),
    .QN(_2188_));
 DFF_X1 _5320_ (.D(_0667_),
    .CK(clknet_leaf_20_pclk),
    .Q(\mem[25] [25]),
    .QN(_2187_));
 DFF_X1 _5321_ (.D(_0668_),
    .CK(clknet_leaf_8_pclk),
    .Q(\mem[25] [26]),
    .QN(_2186_));
 DFF_X1 _5322_ (.D(_0669_),
    .CK(clknet_leaf_0_pclk),
    .Q(\mem[25] [27]),
    .QN(_2185_));
 DFF_X1 _5323_ (.D(_0670_),
    .CK(clknet_leaf_23_pclk),
    .Q(\mem[25] [28]),
    .QN(_2184_));
 DFF_X1 _5324_ (.D(_0671_),
    .CK(clknet_leaf_32_pclk),
    .Q(\mem[25] [29]),
    .QN(_2183_));
 DFF_X1 _5325_ (.D(_0672_),
    .CK(clknet_leaf_19_pclk),
    .Q(\mem[25] [30]),
    .QN(_2182_));
 DFF_X1 _5326_ (.D(_0673_),
    .CK(clknet_leaf_31_pclk),
    .Q(\mem[25] [31]),
    .QN(_2181_));
 DFF_X1 _5327_ (.D(_0674_),
    .CK(clknet_leaf_20_pclk),
    .Q(\mem[7] [0]),
    .QN(_2180_));
 DFF_X1 _5328_ (.D(_0675_),
    .CK(clknet_leaf_27_pclk),
    .Q(\mem[7] [1]),
    .QN(_2179_));
 DFF_X1 _5329_ (.D(_0676_),
    .CK(clknet_leaf_3_pclk),
    .Q(\mem[7] [2]),
    .QN(_2178_));
 DFF_X1 _5330_ (.D(_0677_),
    .CK(clknet_leaf_14_pclk),
    .Q(\mem[7] [3]),
    .QN(_2177_));
 DFF_X1 _5331_ (.D(_0678_),
    .CK(clknet_leaf_21_pclk),
    .Q(\mem[7] [4]),
    .QN(_2176_));
 DFF_X1 _5332_ (.D(_0679_),
    .CK(clknet_leaf_10_pclk),
    .Q(\mem[7] [5]),
    .QN(_2175_));
 DFF_X1 _5333_ (.D(_0680_),
    .CK(clknet_leaf_2_pclk),
    .Q(\mem[7] [6]),
    .QN(_2174_));
 DFF_X1 _5334_ (.D(_0681_),
    .CK(clknet_leaf_27_pclk),
    .Q(\mem[7] [7]),
    .QN(_2173_));
 DFF_X1 _5335_ (.D(_0682_),
    .CK(clknet_leaf_34_pclk),
    .Q(\mem[7] [8]),
    .QN(_2172_));
 DFF_X1 _5336_ (.D(_0683_),
    .CK(clknet_leaf_5_pclk),
    .Q(\mem[7] [9]),
    .QN(_2171_));
 DFF_X1 _5337_ (.D(_0684_),
    .CK(clknet_leaf_17_pclk),
    .Q(\mem[7] [10]),
    .QN(_2170_));
 DFF_X1 _5338_ (.D(_0685_),
    .CK(clknet_leaf_4_pclk),
    .Q(\mem[7] [11]),
    .QN(_2169_));
 DFF_X1 _5339_ (.D(_0686_),
    .CK(clknet_leaf_3_pclk),
    .Q(\mem[7] [12]),
    .QN(_2168_));
 DFF_X1 _5340_ (.D(_0687_),
    .CK(clknet_leaf_29_pclk),
    .Q(\mem[7] [13]),
    .QN(_2167_));
 DFF_X1 _5341_ (.D(_0688_),
    .CK(clknet_leaf_24_pclk),
    .Q(\mem[7] [14]),
    .QN(_2166_));
 DFF_X1 _5342_ (.D(_0689_),
    .CK(clknet_leaf_24_pclk),
    .Q(\mem[7] [15]),
    .QN(_2165_));
 DFF_X1 _5343_ (.D(_0690_),
    .CK(clknet_leaf_12_pclk),
    .Q(\mem[7] [16]),
    .QN(_2164_));
 DFF_X1 _5344_ (.D(_0691_),
    .CK(clknet_leaf_12_pclk),
    .Q(\mem[7] [17]),
    .QN(_2163_));
 DFF_X1 _5345_ (.D(_0692_),
    .CK(clknet_leaf_11_pclk),
    .Q(\mem[7] [18]),
    .QN(_2162_));
 DFF_X1 _5346_ (.D(_0693_),
    .CK(clknet_leaf_4_pclk),
    .Q(\mem[7] [19]),
    .QN(_2161_));
 DFF_X1 _5347_ (.D(_0694_),
    .CK(clknet_leaf_33_pclk),
    .Q(\mem[7] [20]),
    .QN(_2160_));
 DFF_X1 _5348_ (.D(_0695_),
    .CK(clknet_leaf_15_pclk),
    .Q(\mem[7] [21]),
    .QN(_2159_));
 DFF_X1 _5349_ (.D(_0696_),
    .CK(clknet_leaf_9_pclk),
    .Q(\mem[7] [22]),
    .QN(_2158_));
 DFF_X1 _5350_ (.D(_0697_),
    .CK(clknet_leaf_29_pclk),
    .Q(\mem[7] [23]),
    .QN(_2157_));
 DFF_X1 _5351_ (.D(_0698_),
    .CK(clknet_leaf_16_pclk),
    .Q(\mem[7] [24]),
    .QN(_2156_));
 DFF_X1 _5352_ (.D(_0699_),
    .CK(clknet_leaf_12_pclk),
    .Q(\mem[7] [25]),
    .QN(_2155_));
 DFF_X1 _5353_ (.D(_0700_),
    .CK(clknet_leaf_8_pclk),
    .Q(\mem[7] [26]),
    .QN(_2154_));
 DFF_X1 _5354_ (.D(_0701_),
    .CK(clknet_leaf_0_pclk),
    .Q(\mem[7] [27]),
    .QN(_2153_));
 DFF_X1 _5355_ (.D(_0702_),
    .CK(clknet_leaf_24_pclk),
    .Q(\mem[7] [28]),
    .QN(_2152_));
 DFF_X1 _5356_ (.D(_0703_),
    .CK(clknet_leaf_31_pclk),
    .Q(\mem[7] [29]),
    .QN(_2151_));
 DFF_X1 _5357_ (.D(_0704_),
    .CK(clknet_leaf_19_pclk),
    .Q(\mem[7] [30]),
    .QN(_2150_));
 DFF_X1 _5358_ (.D(_0705_),
    .CK(clknet_leaf_31_pclk),
    .Q(\mem[7] [31]),
    .QN(_2149_));
 DFF_X1 _5359_ (.D(_0706_),
    .CK(clknet_leaf_19_pclk),
    .Q(\mem[10] [0]),
    .QN(_2148_));
 DFF_X1 _5360_ (.D(_0707_),
    .CK(clknet_leaf_27_pclk),
    .Q(\mem[10] [1]),
    .QN(_2147_));
 DFF_X1 _5361_ (.D(_0708_),
    .CK(clknet_leaf_3_pclk),
    .Q(\mem[10] [2]),
    .QN(_2146_));
 DFF_X1 _5362_ (.D(_0709_),
    .CK(clknet_leaf_14_pclk),
    .Q(\mem[10] [3]),
    .QN(_2145_));
 DFF_X1 _5363_ (.D(_0710_),
    .CK(clknet_leaf_21_pclk),
    .Q(\mem[10] [4]),
    .QN(_2144_));
 DFF_X1 _5364_ (.D(_0711_),
    .CK(clknet_leaf_10_pclk),
    .Q(\mem[10] [5]),
    .QN(_2143_));
 DFF_X1 _5365_ (.D(_0712_),
    .CK(clknet_leaf_2_pclk),
    .Q(\mem[10] [6]),
    .QN(_2142_));
 DFF_X1 _5366_ (.D(_0713_),
    .CK(clknet_leaf_27_pclk),
    .Q(\mem[10] [7]),
    .QN(_2141_));
 DFF_X1 _5367_ (.D(_0714_),
    .CK(clknet_leaf_34_pclk),
    .Q(\mem[10] [8]),
    .QN(_2140_));
 DFF_X1 _5368_ (.D(_0715_),
    .CK(clknet_leaf_5_pclk),
    .Q(\mem[10] [9]),
    .QN(_2139_));
 DFF_X1 _5369_ (.D(_0716_),
    .CK(clknet_leaf_16_pclk),
    .Q(\mem[10] [10]),
    .QN(_2138_));
 DFF_X1 _5370_ (.D(_0717_),
    .CK(clknet_leaf_4_pclk),
    .Q(\mem[10] [11]),
    .QN(_2137_));
 DFF_X1 _5371_ (.D(_0718_),
    .CK(clknet_leaf_2_pclk),
    .Q(\mem[10] [12]),
    .QN(_2136_));
 DFF_X1 _5372_ (.D(_0719_),
    .CK(clknet_leaf_21_pclk),
    .Q(\mem[10] [13]),
    .QN(_2135_));
 DFF_X1 _5373_ (.D(_0720_),
    .CK(clknet_leaf_26_pclk),
    .Q(\mem[10] [14]),
    .QN(_2134_));
 DFF_X1 _5374_ (.D(_0721_),
    .CK(clknet_leaf_24_pclk),
    .Q(\mem[10] [15]),
    .QN(_2133_));
 DFF_X1 _5375_ (.D(_0722_),
    .CK(clknet_leaf_4_pclk),
    .Q(\mem[10] [16]),
    .QN(_2132_));
 DFF_X1 _5376_ (.D(_0723_),
    .CK(clknet_leaf_13_pclk),
    .Q(\mem[10] [17]),
    .QN(_2131_));
 DFF_X1 _5377_ (.D(_0724_),
    .CK(clknet_leaf_9_pclk),
    .Q(\mem[10] [18]),
    .QN(_2130_));
 DFF_X1 _5378_ (.D(_0725_),
    .CK(clknet_leaf_6_pclk),
    .Q(\mem[10] [19]),
    .QN(_2129_));
 DFF_X1 _5379_ (.D(_0726_),
    .CK(clknet_leaf_33_pclk),
    .Q(\mem[10] [20]),
    .QN(_2128_));
 DFF_X1 _5380_ (.D(_0727_),
    .CK(clknet_leaf_13_pclk),
    .Q(\mem[10] [21]),
    .QN(_2127_));
 DFF_X1 _5381_ (.D(_0728_),
    .CK(clknet_leaf_8_pclk),
    .Q(\mem[10] [22]),
    .QN(_2126_));
 DFF_X1 _5382_ (.D(_0729_),
    .CK(clknet_leaf_29_pclk),
    .Q(\mem[10] [23]),
    .QN(_2125_));
 DFF_X1 _5383_ (.D(_0730_),
    .CK(clknet_leaf_16_pclk),
    .Q(\mem[10] [24]),
    .QN(_2124_));
 DFF_X1 _5384_ (.D(_0731_),
    .CK(clknet_leaf_21_pclk),
    .Q(\mem[10] [25]),
    .QN(_2123_));
 DFF_X1 _5385_ (.D(_0732_),
    .CK(clknet_leaf_8_pclk),
    .Q(\mem[10] [26]),
    .QN(_2122_));
 DFF_X1 _5386_ (.D(_0733_),
    .CK(clknet_leaf_0_pclk),
    .Q(\mem[10] [27]),
    .QN(_2121_));
 DFF_X1 _5387_ (.D(_0734_),
    .CK(clknet_leaf_29_pclk),
    .Q(\mem[10] [28]),
    .QN(_2120_));
 DFF_X1 _5388_ (.D(_0735_),
    .CK(clknet_leaf_33_pclk),
    .Q(\mem[10] [29]),
    .QN(_2119_));
 DFF_X1 _5389_ (.D(_0736_),
    .CK(clknet_leaf_19_pclk),
    .Q(\mem[10] [30]),
    .QN(_2118_));
 DFF_X1 _5390_ (.D(_0737_),
    .CK(clknet_leaf_32_pclk),
    .Q(\mem[10] [31]),
    .QN(_2117_));
 DFF_X1 _5391_ (.D(_0738_),
    .CK(clknet_leaf_20_pclk),
    .Q(\mem[29] [0]),
    .QN(_2116_));
 DFF_X1 _5392_ (.D(_0739_),
    .CK(clknet_leaf_27_pclk),
    .Q(\mem[29] [1]),
    .QN(_2115_));
 DFF_X1 _5393_ (.D(_0740_),
    .CK(clknet_leaf_3_pclk),
    .Q(\mem[29] [2]),
    .QN(_2114_));
 DFF_X1 _5394_ (.D(_0741_),
    .CK(clknet_leaf_15_pclk),
    .Q(\mem[29] [3]),
    .QN(_2113_));
 DFF_X1 _5395_ (.D(_0742_),
    .CK(clknet_leaf_22_pclk),
    .Q(\mem[29] [4]),
    .QN(_2112_));
 DFF_X1 _5396_ (.D(_0743_),
    .CK(clknet_leaf_10_pclk),
    .Q(\mem[29] [5]),
    .QN(_2111_));
 DFF_X1 _5397_ (.D(_0744_),
    .CK(clknet_leaf_1_pclk),
    .Q(\mem[29] [6]),
    .QN(_2110_));
 DFF_X1 _5398_ (.D(_0745_),
    .CK(clknet_leaf_27_pclk),
    .Q(\mem[29] [7]),
    .QN(_2109_));
 DFF_X1 _5399_ (.D(_0746_),
    .CK(clknet_leaf_35_pclk),
    .Q(\mem[29] [8]),
    .QN(_2108_));
 DFF_X1 _5400_ (.D(_0747_),
    .CK(clknet_leaf_5_pclk),
    .Q(\mem[29] [9]),
    .QN(_2107_));
 DFF_X1 _5401_ (.D(_0748_),
    .CK(clknet_leaf_17_pclk),
    .Q(\mem[29] [10]),
    .QN(_2106_));
 DFF_X1 _5402_ (.D(_0749_),
    .CK(clknet_leaf_7_pclk),
    .Q(\mem[29] [11]),
    .QN(_2105_));
 DFF_X1 _5403_ (.D(_0750_),
    .CK(clknet_leaf_31_pclk),
    .Q(\mem[29] [12]),
    .QN(_2104_));
 DFF_X1 _5404_ (.D(_0751_),
    .CK(clknet_leaf_22_pclk),
    .Q(\mem[29] [13]),
    .QN(_2103_));
 DFF_X1 _5405_ (.D(_0752_),
    .CK(clknet_leaf_26_pclk),
    .Q(\mem[29] [14]),
    .QN(_2102_));
 DFF_X1 _5406_ (.D(_0753_),
    .CK(clknet_leaf_24_pclk),
    .Q(\mem[29] [15]),
    .QN(_2101_));
 DFF_X1 _5407_ (.D(_0754_),
    .CK(clknet_leaf_11_pclk),
    .Q(\mem[29] [16]),
    .QN(_2100_));
 DFF_X1 _5408_ (.D(_0755_),
    .CK(clknet_leaf_14_pclk),
    .Q(\mem[29] [17]),
    .QN(_2099_));
 DFF_X1 _5409_ (.D(_0756_),
    .CK(clknet_leaf_11_pclk),
    .Q(\mem[29] [18]),
    .QN(_2098_));
 DFF_X1 _5410_ (.D(_0757_),
    .CK(clknet_leaf_6_pclk),
    .Q(\mem[29] [19]),
    .QN(_2097_));
 DFF_X1 _5411_ (.D(_0758_),
    .CK(clknet_leaf_34_pclk),
    .Q(\mem[29] [20]),
    .QN(_2096_));
 DFF_X1 _5412_ (.D(_0759_),
    .CK(clknet_leaf_20_pclk),
    .Q(\mem[29] [21]),
    .QN(_2095_));
 DFF_X1 _5413_ (.D(_0760_),
    .CK(clknet_leaf_7_pclk),
    .Q(\mem[29] [22]),
    .QN(_2094_));
 DFF_X1 _5414_ (.D(_0761_),
    .CK(clknet_leaf_30_pclk),
    .Q(\mem[29] [23]),
    .QN(_2093_));
 DFF_X1 _5415_ (.D(_0762_),
    .CK(clknet_leaf_16_pclk),
    .Q(\mem[29] [24]),
    .QN(_2092_));
 DFF_X1 _5416_ (.D(_0763_),
    .CK(clknet_leaf_20_pclk),
    .Q(\mem[29] [25]),
    .QN(_2091_));
 DFF_X1 _5417_ (.D(_0764_),
    .CK(clknet_leaf_7_pclk),
    .Q(\mem[29] [26]),
    .QN(_2090_));
 DFF_X1 _5418_ (.D(_0765_),
    .CK(clknet_leaf_35_pclk),
    .Q(\mem[29] [27]),
    .QN(_2089_));
 DFF_X1 _5419_ (.D(_0766_),
    .CK(clknet_leaf_29_pclk),
    .Q(\mem[29] [28]),
    .QN(_2088_));
 DFF_X1 _5420_ (.D(_0767_),
    .CK(clknet_leaf_32_pclk),
    .Q(\mem[29] [29]),
    .QN(_2087_));
 DFF_X1 _5421_ (.D(_0768_),
    .CK(clknet_leaf_19_pclk),
    .Q(\mem[29] [30]),
    .QN(_2086_));
 DFF_X1 _5422_ (.D(_0769_),
    .CK(clknet_leaf_32_pclk),
    .Q(\mem[29] [31]),
    .QN(_2085_));
 DFFR_X1 _5423_ (.D(_0770_),
    .RN(prst_n),
    .CK(clknet_leaf_16_pclk),
    .Q(pslverr),
    .QN(_2084_));
 DFF_X1 _5424_ (.D(_0771_),
    .CK(clknet_leaf_19_pclk),
    .Q(\mem[3] [0]),
    .QN(_2083_));
 DFF_X1 _5425_ (.D(_0772_),
    .CK(clknet_leaf_26_pclk),
    .Q(\mem[3] [1]),
    .QN(_2082_));
 DFF_X1 _5426_ (.D(_0773_),
    .CK(clknet_leaf_12_pclk),
    .Q(\mem[3] [2]),
    .QN(_2081_));
 DFF_X1 _5427_ (.D(_0774_),
    .CK(clknet_leaf_14_pclk),
    .Q(\mem[3] [3]),
    .QN(_2080_));
 DFF_X1 _5428_ (.D(_0775_),
    .CK(clknet_leaf_23_pclk),
    .Q(\mem[3] [4]),
    .QN(_2079_));
 DFF_X1 _5429_ (.D(_0776_),
    .CK(clknet_leaf_10_pclk),
    .Q(\mem[3] [5]),
    .QN(_2078_));
 DFF_X1 _5430_ (.D(_0777_),
    .CK(clknet_leaf_2_pclk),
    .Q(\mem[3] [6]),
    .QN(_2077_));
 DFF_X1 _5431_ (.D(_0778_),
    .CK(clknet_leaf_28_pclk),
    .Q(\mem[3] [7]),
    .QN(_2076_));
 DFF_X1 _5432_ (.D(_0779_),
    .CK(clknet_leaf_33_pclk),
    .Q(\mem[3] [8]),
    .QN(_2075_));
 DFF_X1 _5433_ (.D(_0780_),
    .CK(clknet_leaf_5_pclk),
    .Q(\mem[3] [9]),
    .QN(_2074_));
 DFF_X1 _5434_ (.D(_0781_),
    .CK(clknet_leaf_16_pclk),
    .Q(\mem[3] [10]),
    .QN(_2073_));
 DFF_X1 _5435_ (.D(_0782_),
    .CK(clknet_leaf_4_pclk),
    .Q(\mem[3] [11]),
    .QN(_2072_));
 DFF_X1 _5436_ (.D(_0783_),
    .CK(clknet_leaf_31_pclk),
    .Q(\mem[3] [12]),
    .QN(_2071_));
 DFF_X1 _5437_ (.D(_0784_),
    .CK(clknet_leaf_29_pclk),
    .Q(\mem[3] [13]),
    .QN(_2070_));
 DFF_X1 _5438_ (.D(_0785_),
    .CK(clknet_leaf_25_pclk),
    .Q(\mem[3] [14]),
    .QN(_2069_));
 DFF_X1 _5439_ (.D(_0786_),
    .CK(clknet_leaf_24_pclk),
    .Q(\mem[3] [15]),
    .QN(_2068_));
 DFF_X1 _5440_ (.D(_0787_),
    .CK(clknet_leaf_12_pclk),
    .Q(\mem[3] [16]),
    .QN(_2067_));
 DFF_X1 _5441_ (.D(_0788_),
    .CK(clknet_leaf_13_pclk),
    .Q(\mem[3] [17]),
    .QN(_2066_));
 DFF_X1 _5442_ (.D(_0789_),
    .CK(clknet_leaf_9_pclk),
    .Q(\mem[3] [18]),
    .QN(_2065_));
 DFF_X1 _5443_ (.D(_0790_),
    .CK(clknet_leaf_4_pclk),
    .Q(\mem[3] [19]),
    .QN(_2064_));
 DFF_X1 _5444_ (.D(_0791_),
    .CK(clknet_leaf_33_pclk),
    .Q(\mem[3] [20]),
    .QN(_2063_));
 DFF_X1 _5445_ (.D(_0792_),
    .CK(clknet_leaf_15_pclk),
    .Q(\mem[3] [21]),
    .QN(_2062_));
 DFF_X1 _5446_ (.D(_0793_),
    .CK(clknet_leaf_8_pclk),
    .Q(\mem[3] [22]),
    .QN(_2061_));
 DFF_X1 _5447_ (.D(_0794_),
    .CK(clknet_leaf_30_pclk),
    .Q(\mem[3] [23]),
    .QN(_2060_));
 DFF_X1 _5448_ (.D(_0795_),
    .CK(clknet_leaf_16_pclk),
    .Q(\mem[3] [24]),
    .QN(_2059_));
 DFF_X1 _5449_ (.D(_0796_),
    .CK(clknet_leaf_20_pclk),
    .Q(\mem[3] [25]),
    .QN(_2058_));
 DFF_X1 _5450_ (.D(_0797_),
    .CK(clknet_leaf_9_pclk),
    .Q(\mem[3] [26]),
    .QN(_2057_));
 DFF_X1 _5451_ (.D(_0798_),
    .CK(clknet_leaf_0_pclk),
    .Q(\mem[3] [27]),
    .QN(_2056_));
 DFF_X1 _5452_ (.D(_0799_),
    .CK(clknet_leaf_23_pclk),
    .Q(\mem[3] [28]),
    .QN(_2055_));
 DFF_X1 _5453_ (.D(_0800_),
    .CK(clknet_leaf_33_pclk),
    .Q(\mem[3] [29]),
    .QN(_2054_));
 DFF_X1 _5454_ (.D(_0801_),
    .CK(clknet_leaf_19_pclk),
    .Q(\mem[3] [30]),
    .QN(_2053_));
 DFF_X1 _5455_ (.D(_0802_),
    .CK(clknet_leaf_31_pclk),
    .Q(\mem[3] [31]),
    .QN(_2052_));
 DFF_X1 _5456_ (.D(_0803_),
    .CK(clknet_leaf_18_pclk),
    .Q(\mem[8] [0]),
    .QN(_2051_));
 DFF_X1 _5457_ (.D(_0804_),
    .CK(clknet_leaf_26_pclk),
    .Q(\mem[8] [1]),
    .QN(_2050_));
 DFF_X1 _5458_ (.D(_0805_),
    .CK(clknet_leaf_12_pclk),
    .Q(\mem[8] [2]),
    .QN(_2049_));
 DFF_X1 _5459_ (.D(_0806_),
    .CK(clknet_leaf_15_pclk),
    .Q(\mem[8] [3]),
    .QN(_2048_));
 DFF_X1 _5460_ (.D(_0807_),
    .CK(clknet_leaf_21_pclk),
    .Q(\mem[8] [4]),
    .QN(_2047_));
 DFF_X1 _5461_ (.D(_0808_),
    .CK(clknet_leaf_10_pclk),
    .Q(\mem[8] [5]),
    .QN(_2046_));
 DFF_X1 _5462_ (.D(_0809_),
    .CK(clknet_leaf_2_pclk),
    .Q(\mem[8] [6]),
    .QN(_2045_));
 DFF_X1 _5463_ (.D(_0810_),
    .CK(clknet_leaf_27_pclk),
    .Q(\mem[8] [7]),
    .QN(_2044_));
 DFF_X1 _5464_ (.D(_0811_),
    .CK(clknet_leaf_34_pclk),
    .Q(\mem[8] [8]),
    .QN(_2043_));
 DFF_X1 _5465_ (.D(_0812_),
    .CK(clknet_leaf_2_pclk),
    .Q(\mem[8] [9]),
    .QN(_2042_));
 DFF_X1 _5466_ (.D(_0813_),
    .CK(clknet_leaf_17_pclk),
    .Q(\mem[8] [10]),
    .QN(_2041_));
 DFF_X1 _5467_ (.D(_0814_),
    .CK(clknet_leaf_5_pclk),
    .Q(\mem[8] [11]),
    .QN(_2040_));
 DFF_X1 _5468_ (.D(_0815_),
    .CK(clknet_leaf_30_pclk),
    .Q(\mem[8] [12]),
    .QN(_2039_));
 DFF_X1 _5469_ (.D(_0816_),
    .CK(clknet_leaf_29_pclk),
    .Q(\mem[8] [13]),
    .QN(_2038_));
 DFF_X1 _5470_ (.D(_0817_),
    .CK(clknet_leaf_26_pclk),
    .Q(\mem[8] [14]),
    .QN(_2037_));
 DFF_X1 _5471_ (.D(_0818_),
    .CK(clknet_leaf_24_pclk),
    .Q(\mem[8] [15]),
    .QN(_2036_));
 DFF_X1 _5472_ (.D(_0819_),
    .CK(clknet_leaf_4_pclk),
    .Q(\mem[8] [16]),
    .QN(_2035_));
 DFF_X1 _5473_ (.D(_0820_),
    .CK(clknet_leaf_13_pclk),
    .Q(\mem[8] [17]),
    .QN(_2034_));
 DFF_X1 _5474_ (.D(_0821_),
    .CK(clknet_leaf_9_pclk),
    .Q(\mem[8] [18]),
    .QN(_2033_));
 DFF_X1 _5475_ (.D(_0822_),
    .CK(clknet_leaf_6_pclk),
    .Q(\mem[8] [19]),
    .QN(_2032_));
 DFF_X1 _5476_ (.D(_0823_),
    .CK(clknet_leaf_33_pclk),
    .Q(\mem[8] [20]),
    .QN(_2031_));
 DFF_X1 _5477_ (.D(_0824_),
    .CK(clknet_leaf_13_pclk),
    .Q(\mem[8] [21]),
    .QN(_2030_));
 DFF_X1 _5478_ (.D(_0825_),
    .CK(clknet_leaf_7_pclk),
    .Q(\mem[8] [22]),
    .QN(_2029_));
 DFF_X1 _5479_ (.D(_0826_),
    .CK(clknet_leaf_30_pclk),
    .Q(\mem[8] [23]),
    .QN(_2028_));
 DFF_X1 _5480_ (.D(_0827_),
    .CK(clknet_leaf_16_pclk),
    .Q(\mem[8] [24]),
    .QN(_2027_));
 DFF_X1 _5481_ (.D(_0828_),
    .CK(clknet_leaf_20_pclk),
    .Q(\mem[8] [25]),
    .QN(_2026_));
 DFF_X1 _5482_ (.D(_0829_),
    .CK(clknet_leaf_8_pclk),
    .Q(\mem[8] [26]),
    .QN(_2025_));
 DFF_X1 _5483_ (.D(_0830_),
    .CK(clknet_leaf_35_pclk),
    .Q(\mem[8] [27]),
    .QN(_2024_));
 DFF_X1 _5484_ (.D(_0831_),
    .CK(clknet_leaf_24_pclk),
    .Q(\mem[8] [28]),
    .QN(_2023_));
 DFF_X1 _5485_ (.D(_0832_),
    .CK(clknet_leaf_32_pclk),
    .Q(\mem[8] [29]),
    .QN(_2022_));
 DFF_X1 _5486_ (.D(_0833_),
    .CK(clknet_leaf_19_pclk),
    .Q(\mem[8] [30]),
    .QN(_2021_));
 DFF_X1 _5487_ (.D(_0834_),
    .CK(clknet_leaf_32_pclk),
    .Q(\mem[8] [31]),
    .QN(_2020_));
 DFF_X1 _5488_ (.D(_0835_),
    .CK(clknet_leaf_18_pclk),
    .Q(\mem[5] [0]),
    .QN(_2019_));
 DFF_X1 _5489_ (.D(_0836_),
    .CK(clknet_leaf_26_pclk),
    .Q(\mem[5] [1]),
    .QN(_2018_));
 DFF_X1 _5490_ (.D(_0837_),
    .CK(clknet_leaf_3_pclk),
    .Q(\mem[5] [2]),
    .QN(_2017_));
 DFF_X1 _5491_ (.D(_0838_),
    .CK(clknet_leaf_14_pclk),
    .Q(\mem[5] [3]),
    .QN(_2016_));
 DFF_X1 _5492_ (.D(_0839_),
    .CK(clknet_leaf_22_pclk),
    .Q(\mem[5] [4]),
    .QN(_2015_));
 DFF_X1 _5493_ (.D(_0840_),
    .CK(clknet_leaf_10_pclk),
    .Q(\mem[5] [5]),
    .QN(_2014_));
 DFF_X1 _5494_ (.D(_0841_),
    .CK(clknet_leaf_0_pclk),
    .Q(\mem[5] [6]),
    .QN(_2013_));
 DFF_X1 _5495_ (.D(_0842_),
    .CK(clknet_leaf_29_pclk),
    .Q(\mem[5] [7]),
    .QN(_2012_));
 DFF_X1 _5496_ (.D(_0843_),
    .CK(clknet_leaf_0_pclk),
    .Q(\mem[5] [8]),
    .QN(_2011_));
 DFF_X1 _5497_ (.D(_0844_),
    .CK(clknet_leaf_5_pclk),
    .Q(\mem[5] [9]),
    .QN(_2010_));
 DFF_X1 _5498_ (.D(_0845_),
    .CK(clknet_leaf_17_pclk),
    .Q(\mem[5] [10]),
    .QN(_2009_));
 DFF_X1 _5499_ (.D(_0846_),
    .CK(clknet_leaf_5_pclk),
    .Q(\mem[5] [11]),
    .QN(_2008_));
 DFF_X1 _5500_ (.D(_0847_),
    .CK(clknet_leaf_2_pclk),
    .Q(\mem[5] [12]),
    .QN(_2007_));
 DFF_X1 _5501_ (.D(_0848_),
    .CK(clknet_leaf_29_pclk),
    .Q(\mem[5] [13]),
    .QN(_2006_));
 DFF_X1 _5502_ (.D(_0849_),
    .CK(clknet_leaf_25_pclk),
    .Q(\mem[5] [14]),
    .QN(_2005_));
 DFF_X1 _5503_ (.D(_0850_),
    .CK(clknet_leaf_25_pclk),
    .Q(\mem[5] [15]),
    .QN(_2004_));
 DFF_X1 _5504_ (.D(_0851_),
    .CK(clknet_leaf_11_pclk),
    .Q(\mem[5] [16]),
    .QN(_2003_));
 DFF_X1 _5505_ (.D(_0852_),
    .CK(clknet_leaf_10_pclk),
    .Q(\mem[5] [17]),
    .QN(_2002_));
 DFF_X1 _5506_ (.D(_0853_),
    .CK(clknet_leaf_8_pclk),
    .Q(\mem[5] [18]),
    .QN(_2001_));
 DFF_X1 _5507_ (.D(_0854_),
    .CK(clknet_leaf_5_pclk),
    .Q(\mem[5] [19]),
    .QN(_2000_));
 DFF_X1 _5508_ (.D(_0855_),
    .CK(clknet_leaf_33_pclk),
    .Q(\mem[5] [20]),
    .QN(_1999_));
 DFF_X1 _5509_ (.D(_0856_),
    .CK(clknet_leaf_15_pclk),
    .Q(\mem[5] [21]),
    .QN(_1998_));
 DFF_X1 _5510_ (.D(_0857_),
    .CK(clknet_leaf_7_pclk),
    .Q(\mem[5] [22]),
    .QN(_1997_));
 DFF_X1 _5511_ (.D(_0858_),
    .CK(clknet_leaf_30_pclk),
    .Q(\mem[5] [23]),
    .QN(_1996_));
 DFF_X1 _5512_ (.D(_0859_),
    .CK(clknet_leaf_16_pclk),
    .Q(\mem[5] [24]),
    .QN(_1995_));
 DFF_X1 _5513_ (.D(_0860_),
    .CK(clknet_leaf_12_pclk),
    .Q(\mem[5] [25]),
    .QN(_1994_));
 DFF_X1 _5514_ (.D(_0861_),
    .CK(clknet_leaf_8_pclk),
    .Q(\mem[5] [26]),
    .QN(_1993_));
 DFF_X1 _5515_ (.D(_0862_),
    .CK(clknet_leaf_0_pclk),
    .Q(\mem[5] [27]),
    .QN(_1992_));
 DFF_X1 _5516_ (.D(_0863_),
    .CK(clknet_leaf_24_pclk),
    .Q(\mem[5] [28]),
    .QN(_1991_));
 DFF_X1 _5517_ (.D(_0864_),
    .CK(clknet_leaf_31_pclk),
    .Q(\mem[5] [29]),
    .QN(_1990_));
 DFF_X1 _5518_ (.D(_0865_),
    .CK(clknet_leaf_19_pclk),
    .Q(\mem[5] [30]),
    .QN(_1989_));
 DFF_X1 _5519_ (.D(_0866_),
    .CK(clknet_leaf_31_pclk),
    .Q(\mem[5] [31]),
    .QN(_1988_));
 DFF_X1 _5520_ (.D(_0867_),
    .CK(clknet_leaf_19_pclk),
    .Q(\mem[0] [0]),
    .QN(_1987_));
 DFF_X1 _5521_ (.D(_0868_),
    .CK(clknet_leaf_26_pclk),
    .Q(\mem[0] [1]),
    .QN(_1986_));
 DFF_X1 _5522_ (.D(_0869_),
    .CK(clknet_leaf_30_pclk),
    .Q(\mem[0] [2]),
    .QN(_1985_));
 DFF_X1 _5523_ (.D(_0870_),
    .CK(clknet_leaf_14_pclk),
    .Q(\mem[0] [3]),
    .QN(_1984_));
 DFF_X1 _5524_ (.D(_0871_),
    .CK(clknet_leaf_21_pclk),
    .Q(\mem[0] [4]),
    .QN(_1983_));
 DFF_X1 _5525_ (.D(_0872_),
    .CK(clknet_leaf_10_pclk),
    .Q(\mem[0] [5]),
    .QN(_1982_));
 DFF_X1 _5526_ (.D(_0873_),
    .CK(clknet_leaf_2_pclk),
    .Q(\mem[0] [6]),
    .QN(_1981_));
 DFF_X1 _5527_ (.D(_0874_),
    .CK(clknet_leaf_28_pclk),
    .Q(\mem[0] [7]),
    .QN(_1980_));
 DFF_X1 _5528_ (.D(_0875_),
    .CK(clknet_leaf_33_pclk),
    .Q(\mem[0] [8]),
    .QN(_1979_));
 DFF_X1 _5529_ (.D(_0876_),
    .CK(clknet_leaf_5_pclk),
    .Q(\mem[0] [9]),
    .QN(_1978_));
 DFF_X1 _5530_ (.D(_0877_),
    .CK(clknet_leaf_17_pclk),
    .Q(\mem[0] [10]),
    .QN(_1977_));
 DFF_X1 _5531_ (.D(_0878_),
    .CK(clknet_leaf_4_pclk),
    .Q(\mem[0] [11]),
    .QN(_1976_));
 DFF_X1 _5532_ (.D(_0879_),
    .CK(clknet_leaf_3_pclk),
    .Q(\mem[0] [12]),
    .QN(_1975_));
 DFF_X1 _5533_ (.D(_0880_),
    .CK(clknet_leaf_21_pclk),
    .Q(\mem[0] [13]),
    .QN(_1974_));
 DFF_X1 _5534_ (.D(_0881_),
    .CK(clknet_leaf_25_pclk),
    .Q(\mem[0] [14]),
    .QN(_1973_));
 DFF_X1 _5535_ (.D(_0882_),
    .CK(clknet_leaf_24_pclk),
    .Q(\mem[0] [15]),
    .QN(_1972_));
 DFF_X1 _5536_ (.D(_0883_),
    .CK(clknet_leaf_12_pclk),
    .Q(\mem[0] [16]),
    .QN(_1971_));
 DFF_X1 _5537_ (.D(_0884_),
    .CK(clknet_leaf_10_pclk),
    .Q(\mem[0] [17]),
    .QN(_1970_));
 DFF_X1 _5538_ (.D(_0885_),
    .CK(clknet_leaf_11_pclk),
    .Q(\mem[0] [18]),
    .QN(_1969_));
 DFF_X1 _5539_ (.D(_0886_),
    .CK(clknet_leaf_5_pclk),
    .Q(\mem[0] [19]),
    .QN(_1968_));
 DFF_X1 _5540_ (.D(_0887_),
    .CK(clknet_leaf_33_pclk),
    .Q(\mem[0] [20]),
    .QN(_1967_));
 DFF_X1 _5541_ (.D(_0888_),
    .CK(clknet_leaf_15_pclk),
    .Q(\mem[0] [21]),
    .QN(_1966_));
 DFF_X1 _5542_ (.D(_0889_),
    .CK(clknet_leaf_8_pclk),
    .Q(\mem[0] [22]),
    .QN(_1965_));
 DFF_X1 _5543_ (.D(_0890_),
    .CK(clknet_leaf_29_pclk),
    .Q(\mem[0] [23]),
    .QN(_1964_));
 DFF_X1 _5544_ (.D(_0891_),
    .CK(clknet_leaf_17_pclk),
    .Q(\mem[0] [24]),
    .QN(_1963_));
 DFF_X1 _5545_ (.D(_0892_),
    .CK(clknet_leaf_13_pclk),
    .Q(\mem[0] [25]),
    .QN(_1962_));
 DFF_X1 _5546_ (.D(_0893_),
    .CK(clknet_leaf_8_pclk),
    .Q(\mem[0] [26]),
    .QN(_1961_));
 DFF_X1 _5547_ (.D(_0894_),
    .CK(clknet_leaf_0_pclk),
    .Q(\mem[0] [27]),
    .QN(_1960_));
 DFF_X1 _5548_ (.D(_0895_),
    .CK(clknet_leaf_24_pclk),
    .Q(\mem[0] [28]),
    .QN(_1959_));
 DFF_X1 _5549_ (.D(_0896_),
    .CK(clknet_leaf_33_pclk),
    .Q(\mem[0] [29]),
    .QN(_1958_));
 DFF_X1 _5550_ (.D(_0897_),
    .CK(clknet_leaf_22_pclk),
    .Q(\mem[0] [30]),
    .QN(_1957_));
 DFF_X1 _5551_ (.D(_0898_),
    .CK(clknet_leaf_31_pclk),
    .Q(\mem[0] [31]),
    .QN(_1956_));
 DFF_X1 _5552_ (.D(_0899_),
    .CK(clknet_leaf_20_pclk),
    .Q(\mem[4] [0]),
    .QN(_1955_));
 DFF_X1 _5553_ (.D(_0900_),
    .CK(clknet_leaf_27_pclk),
    .Q(\mem[4] [1]),
    .QN(_1954_));
 DFF_X1 _5554_ (.D(_0901_),
    .CK(clknet_leaf_12_pclk),
    .Q(\mem[4] [2]),
    .QN(_1953_));
 DFF_X1 _5555_ (.D(_0902_),
    .CK(clknet_leaf_14_pclk),
    .Q(\mem[4] [3]),
    .QN(_1952_));
 DFF_X1 _5556_ (.D(_0903_),
    .CK(clknet_leaf_23_pclk),
    .Q(\mem[4] [4]),
    .QN(_1951_));
 DFF_X1 _5557_ (.D(_0904_),
    .CK(clknet_leaf_14_pclk),
    .Q(\mem[4] [5]),
    .QN(_1950_));
 DFF_X1 _5558_ (.D(_0905_),
    .CK(clknet_leaf_2_pclk),
    .Q(\mem[4] [6]),
    .QN(_1949_));
 DFF_X1 _5559_ (.D(_0906_),
    .CK(clknet_leaf_27_pclk),
    .Q(\mem[4] [7]),
    .QN(_1948_));
 DFF_X1 _5560_ (.D(_0907_),
    .CK(clknet_leaf_33_pclk),
    .Q(\mem[4] [8]),
    .QN(_1947_));
 DFF_X1 _5561_ (.D(_0908_),
    .CK(clknet_leaf_4_pclk),
    .Q(\mem[4] [9]),
    .QN(_1946_));
 DFF_X1 _5562_ (.D(_0909_),
    .CK(clknet_leaf_17_pclk),
    .Q(\mem[4] [10]),
    .QN(_1945_));
 DFF_X1 _5563_ (.D(_0910_),
    .CK(clknet_leaf_4_pclk),
    .Q(\mem[4] [11]),
    .QN(_1944_));
 DFF_X1 _5564_ (.D(_0911_),
    .CK(clknet_leaf_3_pclk),
    .Q(\mem[4] [12]),
    .QN(_1943_));
 DFF_X1 _5565_ (.D(_0912_),
    .CK(clknet_leaf_29_pclk),
    .Q(\mem[4] [13]),
    .QN(_1942_));
 DFF_X1 _5566_ (.D(_0913_),
    .CK(clknet_leaf_25_pclk),
    .Q(\mem[4] [14]),
    .QN(_1941_));
 DFF_X1 _5567_ (.D(_0914_),
    .CK(clknet_leaf_24_pclk),
    .Q(\mem[4] [15]),
    .QN(_1940_));
 DFF_X1 _5568_ (.D(_0915_),
    .CK(clknet_leaf_12_pclk),
    .Q(\mem[4] [16]),
    .QN(_1939_));
 DFF_X1 _5569_ (.D(_0916_),
    .CK(clknet_leaf_12_pclk),
    .Q(\mem[4] [17]),
    .QN(_1938_));
 DFF_X1 _5570_ (.D(_0917_),
    .CK(clknet_leaf_9_pclk),
    .Q(\mem[4] [18]),
    .QN(_1937_));
 DFF_X1 _5571_ (.D(_0918_),
    .CK(clknet_leaf_4_pclk),
    .Q(\mem[4] [19]),
    .QN(_1936_));
 DFF_X1 _5572_ (.D(_0919_),
    .CK(clknet_leaf_33_pclk),
    .Q(\mem[4] [20]),
    .QN(_1935_));
 DFF_X1 _5573_ (.D(_0920_),
    .CK(clknet_leaf_15_pclk),
    .Q(\mem[4] [21]),
    .QN(_1934_));
 DFF_X1 _5574_ (.D(_0921_),
    .CK(clknet_leaf_9_pclk),
    .Q(\mem[4] [22]),
    .QN(_1933_));
 DFF_X1 _5575_ (.D(_0922_),
    .CK(clknet_leaf_30_pclk),
    .Q(\mem[4] [23]),
    .QN(_1932_));
 DFF_X1 _5576_ (.D(_0923_),
    .CK(clknet_leaf_17_pclk),
    .Q(\mem[4] [24]),
    .QN(_1931_));
 DFF_X1 _5577_ (.D(_0924_),
    .CK(clknet_leaf_13_pclk),
    .Q(\mem[4] [25]),
    .QN(_1930_));
 DFF_X1 _5578_ (.D(_0925_),
    .CK(clknet_leaf_9_pclk),
    .Q(\mem[4] [26]),
    .QN(_1929_));
 DFF_X1 _5579_ (.D(_0926_),
    .CK(clknet_leaf_0_pclk),
    .Q(\mem[4] [27]),
    .QN(_1928_));
 DFF_X1 _5580_ (.D(_0927_),
    .CK(clknet_leaf_23_pclk),
    .Q(\mem[4] [28]),
    .QN(_1927_));
 DFF_X1 _5581_ (.D(_0928_),
    .CK(clknet_leaf_33_pclk),
    .Q(\mem[4] [29]),
    .QN(_1926_));
 DFF_X1 _5582_ (.D(_0929_),
    .CK(clknet_leaf_22_pclk),
    .Q(\mem[4] [30]),
    .QN(_1925_));
 DFF_X1 _5583_ (.D(_0930_),
    .CK(clknet_leaf_32_pclk),
    .Q(\mem[4] [31]),
    .QN(_1924_));
 DFF_X1 _5584_ (.D(_0931_),
    .CK(clknet_leaf_20_pclk),
    .Q(\mem[6] [0]),
    .QN(_1923_));
 DFF_X1 _5585_ (.D(_0932_),
    .CK(clknet_leaf_27_pclk),
    .Q(\mem[6] [1]),
    .QN(_1922_));
 DFF_X1 _5586_ (.D(_0933_),
    .CK(clknet_leaf_3_pclk),
    .Q(\mem[6] [2]),
    .QN(_1921_));
 DFF_X1 _5587_ (.D(_0934_),
    .CK(clknet_leaf_13_pclk),
    .Q(\mem[6] [3]),
    .QN(_1920_));
 DFF_X1 _5588_ (.D(_0935_),
    .CK(clknet_leaf_23_pclk),
    .Q(\mem[6] [4]),
    .QN(_1919_));
 DFF_X1 _5589_ (.D(_0936_),
    .CK(clknet_leaf_10_pclk),
    .Q(\mem[6] [5]),
    .QN(_1918_));
 DFF_X1 _5590_ (.D(_0937_),
    .CK(clknet_leaf_2_pclk),
    .Q(\mem[6] [6]),
    .QN(_1917_));
 DFF_X1 _5591_ (.D(_0938_),
    .CK(clknet_leaf_28_pclk),
    .Q(\mem[6] [7]),
    .QN(_1916_));
 DFF_X1 _5592_ (.D(_0939_),
    .CK(clknet_leaf_0_pclk),
    .Q(\mem[6] [8]),
    .QN(_1915_));
 DFF_X1 _5593_ (.D(_0940_),
    .CK(clknet_leaf_4_pclk),
    .Q(\mem[6] [9]),
    .QN(_1914_));
 DFF_X1 _5594_ (.D(_0941_),
    .CK(clknet_leaf_15_pclk),
    .Q(\mem[6] [10]),
    .QN(_1913_));
 DFF_X1 _5595_ (.D(_0942_),
    .CK(clknet_leaf_4_pclk),
    .Q(\mem[6] [11]),
    .QN(_1912_));
 DFF_X1 _5596_ (.D(_0943_),
    .CK(clknet_leaf_2_pclk),
    .Q(\mem[6] [12]),
    .QN(_1911_));
 DFF_X1 _5597_ (.D(_0944_),
    .CK(clknet_leaf_29_pclk),
    .Q(\mem[6] [13]),
    .QN(_1910_));
 DFF_X1 _5598_ (.D(_0945_),
    .CK(clknet_leaf_25_pclk),
    .Q(\mem[6] [14]),
    .QN(_1909_));
 DFF_X1 _5599_ (.D(_0946_),
    .CK(clknet_leaf_25_pclk),
    .Q(\mem[6] [15]),
    .QN(_1908_));
 DFF_X1 _5600_ (.D(_0947_),
    .CK(clknet_leaf_12_pclk),
    .Q(\mem[6] [16]),
    .QN(_1907_));
 DFF_X1 _5601_ (.D(_0948_),
    .CK(clknet_leaf_12_pclk),
    .Q(\mem[6] [17]),
    .QN(_1906_));
 DFF_X1 _5602_ (.D(_0949_),
    .CK(clknet_leaf_11_pclk),
    .Q(\mem[6] [18]),
    .QN(_1905_));
 DFF_X1 _5603_ (.D(_0950_),
    .CK(clknet_leaf_6_pclk),
    .Q(\mem[6] [19]),
    .QN(_1904_));
 DFF_X1 _5604_ (.D(_0951_),
    .CK(clknet_leaf_33_pclk),
    .Q(\mem[6] [20]),
    .QN(_1903_));
 DFF_X1 _5605_ (.D(_0952_),
    .CK(clknet_leaf_15_pclk),
    .Q(\mem[6] [21]),
    .QN(_1902_));
 DFF_X1 _5606_ (.D(_0953_),
    .CK(clknet_leaf_8_pclk),
    .Q(\mem[6] [22]),
    .QN(_1901_));
 DFF_X1 _5607_ (.D(_0954_),
    .CK(clknet_leaf_29_pclk),
    .Q(\mem[6] [23]),
    .QN(_1900_));
 DFF_X1 _5608_ (.D(_0955_),
    .CK(clknet_leaf_17_pclk),
    .Q(\mem[6] [24]),
    .QN(_1899_));
 DFF_X1 _5609_ (.D(_0956_),
    .CK(clknet_leaf_21_pclk),
    .Q(\mem[6] [25]),
    .QN(_1898_));
 DFF_X1 _5610_ (.D(_0957_),
    .CK(clknet_leaf_9_pclk),
    .Q(\mem[6] [26]),
    .QN(_1897_));
 DFF_X1 _5611_ (.D(_0958_),
    .CK(clknet_leaf_0_pclk),
    .Q(\mem[6] [27]),
    .QN(_1896_));
 DFF_X1 _5612_ (.D(_0959_),
    .CK(clknet_leaf_23_pclk),
    .Q(\mem[6] [28]),
    .QN(_1895_));
 DFF_X1 _5613_ (.D(_0960_),
    .CK(clknet_leaf_31_pclk),
    .Q(\mem[6] [29]),
    .QN(_1894_));
 DFF_X1 _5614_ (.D(_0961_),
    .CK(clknet_leaf_18_pclk),
    .Q(\mem[6] [30]),
    .QN(_1893_));
 DFF_X1 _5615_ (.D(_0962_),
    .CK(clknet_leaf_31_pclk),
    .Q(\mem[6] [31]),
    .QN(_1892_));
 DFF_X1 _5616_ (.D(_0963_),
    .CK(clknet_leaf_18_pclk),
    .Q(\mem[13] [0]),
    .QN(_1891_));
 DFF_X1 _5617_ (.D(_0964_),
    .CK(clknet_leaf_26_pclk),
    .Q(\mem[13] [1]),
    .QN(_1890_));
 DFF_X1 _5618_ (.D(_0965_),
    .CK(clknet_leaf_3_pclk),
    .Q(\mem[13] [2]),
    .QN(_1889_));
 DFF_X1 _5619_ (.D(_0966_),
    .CK(clknet_leaf_14_pclk),
    .Q(\mem[13] [3]),
    .QN(_1888_));
 DFF_X1 _5620_ (.D(_0967_),
    .CK(clknet_leaf_20_pclk),
    .Q(\mem[13] [4]),
    .QN(_1887_));
 DFF_X1 _5621_ (.D(_0968_),
    .CK(clknet_leaf_10_pclk),
    .Q(\mem[13] [5]),
    .QN(_1886_));
 DFF_X1 _5622_ (.D(_0969_),
    .CK(clknet_leaf_1_pclk),
    .Q(\mem[13] [6]),
    .QN(_1885_));
 DFF_X1 _5623_ (.D(_0970_),
    .CK(clknet_leaf_27_pclk),
    .Q(\mem[13] [7]),
    .QN(_1884_));
 DFF_X1 _5624_ (.D(_0971_),
    .CK(clknet_leaf_34_pclk),
    .Q(\mem[13] [8]),
    .QN(_1883_));
 DFF_X1 _5625_ (.D(_0972_),
    .CK(clknet_leaf_1_pclk),
    .Q(\mem[13] [9]),
    .QN(_1882_));
 DFF_X1 _5626_ (.D(_0973_),
    .CK(clknet_leaf_18_pclk),
    .Q(\mem[13] [10]),
    .QN(_1881_));
 DFF_X1 _5627_ (.D(_0974_),
    .CK(clknet_leaf_6_pclk),
    .Q(\mem[13] [11]),
    .QN(_1880_));
 DFF_X1 _5628_ (.D(_0975_),
    .CK(clknet_leaf_30_pclk),
    .Q(\mem[13] [12]),
    .QN(_1879_));
 DFF_X1 _5629_ (.D(_0976_),
    .CK(clknet_leaf_21_pclk),
    .Q(\mem[13] [13]),
    .QN(_1878_));
 DFF_X1 _5630_ (.D(_0977_),
    .CK(clknet_leaf_26_pclk),
    .Q(\mem[13] [14]),
    .QN(_1877_));
 DFF_X1 _5631_ (.D(_0978_),
    .CK(clknet_leaf_25_pclk),
    .Q(\mem[13] [15]),
    .QN(_1876_));
 DFF_X1 _5632_ (.D(_0979_),
    .CK(clknet_leaf_4_pclk),
    .Q(\mem[13] [16]),
    .QN(_1875_));
 DFF_X1 _5633_ (.D(_0980_),
    .CK(clknet_leaf_13_pclk),
    .Q(\mem[13] [17]),
    .QN(_1874_));
 DFF_X1 _5634_ (.D(_0981_),
    .CK(clknet_leaf_9_pclk),
    .Q(\mem[13] [18]),
    .QN(_1873_));
 DFF_X1 _5635_ (.D(_0982_),
    .CK(clknet_leaf_6_pclk),
    .Q(\mem[13] [19]),
    .QN(_1872_));
 DFF_X1 _5636_ (.D(_0983_),
    .CK(clknet_leaf_31_pclk),
    .Q(\mem[13] [20]),
    .QN(_1871_));
 DFF_X1 _5637_ (.D(_0984_),
    .CK(clknet_leaf_13_pclk),
    .Q(\mem[13] [21]),
    .QN(_1870_));
 DFF_X1 _5638_ (.D(_0985_),
    .CK(clknet_leaf_7_pclk),
    .Q(\mem[13] [22]),
    .QN(_1869_));
 DFF_X1 _5639_ (.D(_0986_),
    .CK(clknet_leaf_30_pclk),
    .Q(\mem[13] [23]),
    .QN(_1868_));
 DFF_X1 _5640_ (.D(_0987_),
    .CK(clknet_leaf_16_pclk),
    .Q(\mem[13] [24]),
    .QN(_1867_));
 DFF_X1 _5641_ (.D(_0988_),
    .CK(clknet_leaf_20_pclk),
    .Q(\mem[13] [25]),
    .QN(_1866_));
 DFF_X1 _5642_ (.D(_0989_),
    .CK(clknet_leaf_8_pclk),
    .Q(\mem[13] [26]),
    .QN(_1865_));
 DFF_X1 _5643_ (.D(_0990_),
    .CK(clknet_leaf_0_pclk),
    .Q(\mem[13] [27]),
    .QN(_1864_));
 DFF_X1 _5644_ (.D(_0991_),
    .CK(clknet_leaf_22_pclk),
    .Q(\mem[13] [28]),
    .QN(_1863_));
 DFF_X1 _5645_ (.D(_0992_),
    .CK(clknet_leaf_32_pclk),
    .Q(\mem[13] [29]),
    .QN(_1862_));
 DFF_X1 _5646_ (.D(_0993_),
    .CK(clknet_leaf_19_pclk),
    .Q(\mem[13] [30]),
    .QN(_1861_));
 DFF_X1 _5647_ (.D(_0994_),
    .CK(clknet_leaf_32_pclk),
    .Q(\mem[13] [31]),
    .QN(_1860_));
 DFF_X1 _5648_ (.D(_0995_),
    .CK(clknet_leaf_18_pclk),
    .Q(\mem[14] [0]),
    .QN(_1859_));
 DFF_X1 _5649_ (.D(_0996_),
    .CK(clknet_leaf_25_pclk),
    .Q(\mem[14] [1]),
    .QN(_1858_));
 DFF_X1 _5650_ (.D(_0997_),
    .CK(clknet_leaf_12_pclk),
    .Q(\mem[14] [2]),
    .QN(_1857_));
 DFF_X1 _5651_ (.D(_0998_),
    .CK(clknet_leaf_15_pclk),
    .Q(\mem[14] [3]),
    .QN(_1856_));
 DFF_X1 _5652_ (.D(_0999_),
    .CK(clknet_leaf_22_pclk),
    .Q(\mem[14] [4]),
    .QN(_1855_));
 DFF_X1 _5653_ (.D(_1000_),
    .CK(clknet_leaf_9_pclk),
    .Q(\mem[14] [5]),
    .QN(_1854_));
 DFF_X1 _5654_ (.D(_1001_),
    .CK(clknet_leaf_2_pclk),
    .Q(\mem[14] [6]),
    .QN(_1853_));
 DFF_X1 _5655_ (.D(_1002_),
    .CK(clknet_leaf_27_pclk),
    .Q(\mem[14] [7]),
    .QN(_1852_));
 DFF_X1 _5656_ (.D(_1003_),
    .CK(clknet_leaf_34_pclk),
    .Q(\mem[14] [8]),
    .QN(_1851_));
 DFF_X1 _5657_ (.D(_1004_),
    .CK(clknet_leaf_1_pclk),
    .Q(\mem[14] [9]),
    .QN(_1850_));
 DFF_X1 _5658_ (.D(_1005_),
    .CK(clknet_leaf_17_pclk),
    .Q(\mem[14] [10]),
    .QN(_1849_));
 DFF_X1 _5659_ (.D(_1006_),
    .CK(clknet_leaf_5_pclk),
    .Q(\mem[14] [11]),
    .QN(_1848_));
 DFF_X1 _5660_ (.D(_1007_),
    .CK(clknet_leaf_31_pclk),
    .Q(\mem[14] [12]),
    .QN(_1847_));
 DFF_X1 _5661_ (.D(_1008_),
    .CK(clknet_leaf_22_pclk),
    .Q(\mem[14] [13]),
    .QN(_1846_));
 DFF_X1 _5662_ (.D(_1009_),
    .CK(clknet_leaf_26_pclk),
    .Q(\mem[14] [14]),
    .QN(_1845_));
 DFF_X1 _5663_ (.D(_1010_),
    .CK(clknet_leaf_25_pclk),
    .Q(\mem[14] [15]),
    .QN(_1844_));
 DFF_X1 _5664_ (.D(_1011_),
    .CK(clknet_leaf_3_pclk),
    .Q(\mem[14] [16]),
    .QN(_1843_));
 DFF_X1 _5665_ (.D(_1012_),
    .CK(clknet_leaf_13_pclk),
    .Q(\mem[14] [17]),
    .QN(_1842_));
 DFF_X1 _5666_ (.D(_1013_),
    .CK(clknet_leaf_8_pclk),
    .Q(\mem[14] [18]),
    .QN(_1841_));
 DFF_X1 _5667_ (.D(_1014_),
    .CK(clknet_leaf_6_pclk),
    .Q(\mem[14] [19]),
    .QN(_1840_));
 DFF_X1 _5668_ (.D(_1015_),
    .CK(clknet_leaf_34_pclk),
    .Q(\mem[14] [20]),
    .QN(_1839_));
 DFF_X1 _5669_ (.D(_1016_),
    .CK(clknet_leaf_15_pclk),
    .Q(\mem[14] [21]),
    .QN(_1838_));
 DFF_X1 _5670_ (.D(_1017_),
    .CK(clknet_leaf_7_pclk),
    .Q(\mem[14] [22]),
    .QN(_1837_));
 DFF_X1 _5671_ (.D(_1018_),
    .CK(clknet_leaf_29_pclk),
    .Q(\mem[14] [23]),
    .QN(_1836_));
 DFF_X1 _5672_ (.D(_1019_),
    .CK(clknet_leaf_16_pclk),
    .Q(\mem[14] [24]),
    .QN(_1835_));
 DFF_X1 _5673_ (.D(_1020_),
    .CK(clknet_leaf_20_pclk),
    .Q(\mem[14] [25]),
    .QN(_1834_));
 DFF_X1 _5674_ (.D(_1021_),
    .CK(clknet_leaf_9_pclk),
    .Q(\mem[14] [26]),
    .QN(_1833_));
 DFF_X1 _5675_ (.D(_1022_),
    .CK(clknet_leaf_0_pclk),
    .Q(\mem[14] [27]),
    .QN(_1832_));
 DFF_X1 _5676_ (.D(_1023_),
    .CK(clknet_leaf_24_pclk),
    .Q(\mem[14] [28]),
    .QN(_1831_));
 DFF_X1 _5677_ (.D(_1024_),
    .CK(clknet_leaf_32_pclk),
    .Q(\mem[14] [29]),
    .QN(_1830_));
 DFF_X1 _5678_ (.D(_1025_),
    .CK(clknet_leaf_19_pclk),
    .Q(\mem[14] [30]),
    .QN(_1829_));
 DFF_X1 _5679_ (.D(_1026_),
    .CK(clknet_leaf_32_pclk),
    .Q(\mem[14] [31]),
    .QN(_1828_));
 DFF_X1 _5680_ (.D(_1027_),
    .CK(clknet_leaf_18_pclk),
    .Q(\mem[11] [0]),
    .QN(_1827_));
 DFF_X1 _5681_ (.D(_1028_),
    .CK(clknet_leaf_25_pclk),
    .Q(\mem[11] [1]),
    .QN(_1826_));
 DFF_X1 _5682_ (.D(_1029_),
    .CK(clknet_leaf_12_pclk),
    .Q(\mem[11] [2]),
    .QN(_1825_));
 DFF_X1 _5683_ (.D(_1030_),
    .CK(clknet_leaf_14_pclk),
    .Q(\mem[11] [3]),
    .QN(_1824_));
 DFF_X1 _5684_ (.D(_1031_),
    .CK(clknet_leaf_21_pclk),
    .Q(\mem[11] [4]),
    .QN(_1823_));
 DFF_X1 _5685_ (.D(_1032_),
    .CK(clknet_leaf_14_pclk),
    .Q(\mem[11] [5]),
    .QN(_1822_));
 DFF_X1 _5686_ (.D(_1033_),
    .CK(clknet_leaf_1_pclk),
    .Q(\mem[11] [6]),
    .QN(_1821_));
 DFF_X1 _5687_ (.D(_1034_),
    .CK(clknet_leaf_28_pclk),
    .Q(\mem[11] [7]),
    .QN(_1820_));
 DFF_X1 _5688_ (.D(_1035_),
    .CK(clknet_leaf_35_pclk),
    .Q(\mem[11] [8]),
    .QN(_1819_));
 DFF_X1 _5689_ (.D(_1036_),
    .CK(clknet_leaf_1_pclk),
    .Q(\mem[11] [9]),
    .QN(_1818_));
 DFF_X1 _5690_ (.D(_1037_),
    .CK(clknet_leaf_18_pclk),
    .Q(\mem[11] [10]),
    .QN(_1817_));
 DFF_X1 _5691_ (.D(_1038_),
    .CK(clknet_leaf_4_pclk),
    .Q(\mem[11] [11]),
    .QN(_1816_));
 DFF_X1 _5692_ (.D(_1039_),
    .CK(clknet_leaf_3_pclk),
    .Q(\mem[11] [12]),
    .QN(_1815_));
 DFF_X1 _5693_ (.D(_1040_),
    .CK(clknet_leaf_21_pclk),
    .Q(\mem[11] [13]),
    .QN(_1814_));
 DFF_X1 _5694_ (.D(_1041_),
    .CK(clknet_leaf_25_pclk),
    .Q(\mem[11] [14]),
    .QN(_1813_));
 DFF_X1 _5695_ (.D(_1042_),
    .CK(clknet_leaf_24_pclk),
    .Q(\mem[11] [15]),
    .QN(_1812_));
 DFF_X1 _5696_ (.D(_1043_),
    .CK(clknet_leaf_4_pclk),
    .Q(\mem[11] [16]),
    .QN(_1811_));
 DFF_X1 _5697_ (.D(_1044_),
    .CK(clknet_leaf_10_pclk),
    .Q(\mem[11] [17]),
    .QN(_1810_));
 DFF_X1 _5698_ (.D(_1045_),
    .CK(clknet_leaf_9_pclk),
    .Q(\mem[11] [18]),
    .QN(_1809_));
 DFF_X1 _5699_ (.D(_1046_),
    .CK(clknet_leaf_6_pclk),
    .Q(\mem[11] [19]),
    .QN(_1808_));
 DFF_X1 _5700_ (.D(_1047_),
    .CK(clknet_leaf_0_pclk),
    .Q(\mem[11] [20]),
    .QN(_1807_));
 DFF_X1 _5701_ (.D(_1048_),
    .CK(clknet_leaf_15_pclk),
    .Q(\mem[11] [21]),
    .QN(_1806_));
 DFF_X1 _5702_ (.D(_1049_),
    .CK(clknet_leaf_7_pclk),
    .Q(\mem[11] [22]),
    .QN(_1805_));
 DFF_X1 _5703_ (.D(_1050_),
    .CK(clknet_leaf_29_pclk),
    .Q(\mem[11] [23]),
    .QN(_1804_));
 DFF_X1 _5704_ (.D(_1051_),
    .CK(clknet_leaf_17_pclk),
    .Q(\mem[11] [24]),
    .QN(_1803_));
 DFF_X1 _5705_ (.D(_1052_),
    .CK(clknet_leaf_20_pclk),
    .Q(\mem[11] [25]),
    .QN(_1802_));
 DFF_X1 _5706_ (.D(_1053_),
    .CK(clknet_leaf_7_pclk),
    .Q(\mem[11] [26]),
    .QN(_1801_));
 DFF_X1 _5707_ (.D(_1054_),
    .CK(clknet_leaf_1_pclk),
    .Q(\mem[11] [27]),
    .QN(_1800_));
 DFF_X1 _5708_ (.D(_1055_),
    .CK(clknet_leaf_23_pclk),
    .Q(\mem[11] [28]),
    .QN(_1799_));
 DFF_X1 _5709_ (.D(_1056_),
    .CK(clknet_leaf_32_pclk),
    .Q(\mem[11] [29]),
    .QN(_1798_));
 DFF_X1 _5710_ (.D(_1057_),
    .CK(clknet_leaf_19_pclk),
    .Q(\mem[11] [30]),
    .QN(_1797_));
 DFF_X1 _5711_ (.D(_1058_),
    .CK(clknet_leaf_32_pclk),
    .Q(\mem[11] [31]),
    .QN(_2854_));
 DFFR_X1 _5712_ (.D(next_state[0]),
    .RN(prst_n),
    .CK(clknet_leaf_18_pclk),
    .Q(present_state[0]),
    .QN(_0001_));
 DFFR_X1 _5713_ (.D(next_state[1]),
    .RN(prst_n),
    .CK(clknet_leaf_18_pclk),
    .Q(present_state[1]),
    .QN(_0000_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Right_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Right_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Right_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Right_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Right_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Right_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Right_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Right_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Right_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Right_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Right_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Right_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_Right_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_Right_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_Right_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_Right_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_Right_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_Right_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_Right_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_Right_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_Right_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_Right_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_Right_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_Right_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_Right_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_Right_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_Right_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_Right_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_Right_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_Right_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_Right_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_Right_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_Right_69 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_Right_70 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_Right_71 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_Right_72 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_Right_73 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_Right_74 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_Right_75 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_Right_76 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_Right_77 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_Right_78 ();
 TAPCELL_X1 PHY_EDGE_ROW_79_Right_79 ();
 TAPCELL_X1 PHY_EDGE_ROW_80_Right_80 ();
 TAPCELL_X1 PHY_EDGE_ROW_81_Right_81 ();
 TAPCELL_X1 PHY_EDGE_ROW_82_Right_82 ();
 TAPCELL_X1 PHY_EDGE_ROW_83_Right_83 ();
 TAPCELL_X1 PHY_EDGE_ROW_84_Right_84 ();
 TAPCELL_X1 PHY_EDGE_ROW_85_Right_85 ();
 TAPCELL_X1 PHY_EDGE_ROW_86_Right_86 ();
 TAPCELL_X1 PHY_EDGE_ROW_87_Right_87 ();
 TAPCELL_X1 PHY_EDGE_ROW_88_Right_88 ();
 TAPCELL_X1 PHY_EDGE_ROW_89_Right_89 ();
 TAPCELL_X1 PHY_EDGE_ROW_90_Right_90 ();
 TAPCELL_X1 PHY_EDGE_ROW_91_Right_91 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_92 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_93 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_94 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_95 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_96 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_97 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_98 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_99 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_100 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_101 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_102 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_103 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_104 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_105 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_106 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_107 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_108 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_109 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_110 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_111 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_112 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_113 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_114 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_115 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_116 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_117 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_118 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_119 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_120 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_121 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_122 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_123 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Left_124 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Left_125 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Left_126 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Left_127 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Left_128 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Left_129 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Left_130 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Left_131 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Left_132 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Left_133 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Left_134 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Left_135 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Left_136 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Left_137 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Left_138 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Left_139 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Left_140 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_Left_141 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_Left_142 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_Left_143 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_Left_144 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_Left_145 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_Left_146 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_Left_147 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_Left_148 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_Left_149 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_Left_150 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_Left_151 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_Left_152 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_Left_153 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_Left_154 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_Left_155 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_Left_156 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_Left_157 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_Left_158 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_Left_159 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_Left_160 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_Left_161 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_Left_162 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_Left_163 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_Left_164 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_Left_165 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_Left_166 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_Left_167 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_Left_168 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_Left_169 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_Left_170 ();
 TAPCELL_X1 PHY_EDGE_ROW_79_Left_171 ();
 TAPCELL_X1 PHY_EDGE_ROW_80_Left_172 ();
 TAPCELL_X1 PHY_EDGE_ROW_81_Left_173 ();
 TAPCELL_X1 PHY_EDGE_ROW_82_Left_174 ();
 TAPCELL_X1 PHY_EDGE_ROW_83_Left_175 ();
 TAPCELL_X1 PHY_EDGE_ROW_84_Left_176 ();
 TAPCELL_X1 PHY_EDGE_ROW_85_Left_177 ();
 TAPCELL_X1 PHY_EDGE_ROW_86_Left_178 ();
 TAPCELL_X1 PHY_EDGE_ROW_87_Left_179 ();
 TAPCELL_X1 PHY_EDGE_ROW_88_Left_180 ();
 TAPCELL_X1 PHY_EDGE_ROW_89_Left_181 ();
 TAPCELL_X1 PHY_EDGE_ROW_90_Left_182 ();
 TAPCELL_X1 PHY_EDGE_ROW_91_Left_183 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_184 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_2_185 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_4_186 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_6_187 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_8_188 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_10_189 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_12_190 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_14_191 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_16_192 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_18_193 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_20_194 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_22_195 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_24_196 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_26_197 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_28_198 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_30_199 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_32_200 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_34_201 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_36_202 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_38_203 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_40_204 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_42_205 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_44_206 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_46_207 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_48_208 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_50_209 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_52_210 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_54_211 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_56_212 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_58_213 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_60_214 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_62_215 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_64_216 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_66_217 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_68_218 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_70_219 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_72_220 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_74_221 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_76_222 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_78_223 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_80_224 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_82_225 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_84_226 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_86_227 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_88_228 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_90_229 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_91_230 ();
 BUF_X4 load_slew1 (.A(_1091_),
    .Z(net1));
 BUF_X4 load_slew2 (.A(_1090_),
    .Z(net2));
 BUF_X4 load_slew3 (.A(_1131_),
    .Z(net3));
 BUF_X4 load_slew4 (.A(_1131_),
    .Z(net4));
 BUF_X4 load_slew5 (.A(_1116_),
    .Z(net5));
 BUF_X4 load_slew6 (.A(_1116_),
    .Z(net6));
 BUF_X4 max_cap7 (.A(_1101_),
    .Z(net7));
 BUF_X4 max_cap8 (.A(_1101_),
    .Z(net8));
 BUF_X4 max_cap9 (.A(net10),
    .Z(net9));
 BUF_X4 max_cap10 (.A(net11),
    .Z(net10));
 BUF_X4 load_slew11 (.A(_1099_),
    .Z(net11));
 BUF_X4 max_cap12 (.A(_1093_),
    .Z(net12));
 BUF_X4 max_cap13 (.A(_1093_),
    .Z(net13));
 BUF_X4 max_cap14 (.A(_1077_),
    .Z(net14));
 BUF_X4 load_slew15 (.A(_1077_),
    .Z(net15));
 BUF_X4 load_slew16 (.A(net18),
    .Z(net16));
 BUF_X4 max_cap17 (.A(net18),
    .Z(net17));
 BUF_X4 max_cap18 (.A(_1149_),
    .Z(net18));
 BUF_X4 load_slew19 (.A(net20),
    .Z(net19));
 BUF_X4 max_cap20 (.A(net22),
    .Z(net20));
 BUF_X4 load_slew21 (.A(net22),
    .Z(net21));
 BUF_X4 max_cap22 (.A(_1148_),
    .Z(net22));
 BUF_X4 load_slew23 (.A(net24),
    .Z(net23));
 BUF_X2 wire24 (.A(_1145_),
    .Z(net24));
 BUF_X4 max_cap25 (.A(_1143_),
    .Z(net25));
 BUF_X4 load_slew26 (.A(_1143_),
    .Z(net26));
 BUF_X4 max_cap27 (.A(net28),
    .Z(net27));
 BUF_X4 load_slew28 (.A(_1142_),
    .Z(net28));
 BUF_X4 max_cap29 (.A(net30),
    .Z(net29));
 BUF_X4 max_cap30 (.A(_1142_),
    .Z(net30));
 BUF_X4 load_slew31 (.A(net34),
    .Z(net31));
 BUF_X4 max_cap32 (.A(net34),
    .Z(net32));
 BUF_X4 max_cap33 (.A(_1141_),
    .Z(net33));
 BUF_X4 max_cap34 (.A(_1141_),
    .Z(net34));
 BUF_X4 load_slew35 (.A(_1140_),
    .Z(net35));
 BUF_X2 wire36 (.A(_1140_),
    .Z(net36));
 BUF_X4 load_slew37 (.A(net38),
    .Z(net37));
 BUF_X4 max_cap38 (.A(_1139_),
    .Z(net38));
 BUF_X4 max_cap39 (.A(_1139_),
    .Z(net39));
 BUF_X2 load_slew40 (.A(_1137_),
    .Z(net40));
 BUF_X4 max_cap41 (.A(net42),
    .Z(net41));
 BUF_X4 max_cap42 (.A(_1137_),
    .Z(net42));
 BUF_X4 load_slew43 (.A(_1134_),
    .Z(net43));
 BUF_X4 max_cap44 (.A(_1134_),
    .Z(net44));
 BUF_X4 load_slew45 (.A(_1133_),
    .Z(net45));
 BUF_X4 max_cap46 (.A(_1133_),
    .Z(net46));
 BUF_X4 load_slew47 (.A(_1125_),
    .Z(net47));
 BUF_X4 max_cap48 (.A(net49),
    .Z(net48));
 BUF_X4 load_slew49 (.A(_1125_),
    .Z(net49));
 BUF_X4 max_cap50 (.A(net52),
    .Z(net50));
 BUF_X2 wire51 (.A(net52),
    .Z(net51));
 BUF_X4 load_slew52 (.A(_1120_),
    .Z(net52));
 BUF_X2 wire53 (.A(_1118_),
    .Z(net53));
 BUF_X4 max_cap54 (.A(_1118_),
    .Z(net54));
 BUF_X4 max_cap55 (.A(_1118_),
    .Z(net55));
 BUF_X4 max_cap56 (.A(net57),
    .Z(net56));
 BUF_X2 wire57 (.A(_1113_),
    .Z(net57));
 BUF_X4 max_cap58 (.A(_1113_),
    .Z(net58));
 BUF_X4 load_slew59 (.A(net60),
    .Z(net59));
 BUF_X2 wire60 (.A(_1111_),
    .Z(net60));
 BUF_X4 max_cap61 (.A(net62),
    .Z(net61));
 BUF_X4 load_slew62 (.A(_1109_),
    .Z(net62));
 BUF_X4 max_cap63 (.A(net64),
    .Z(net63));
 BUF_X4 max_cap64 (.A(net65),
    .Z(net64));
 BUF_X4 max_cap65 (.A(_1107_),
    .Z(net65));
 BUF_X4 max_cap66 (.A(_1105_),
    .Z(net66));
 BUF_X4 max_cap67 (.A(_1105_),
    .Z(net67));
 BUF_X4 load_slew68 (.A(net70),
    .Z(net68));
 BUF_X4 max_cap69 (.A(net70),
    .Z(net69));
 BUF_X4 max_cap70 (.A(_1103_),
    .Z(net70));
 BUF_X4 clkbuf_leaf_0_pclk (.A(clknet_2_0__leaf_pclk),
    .Z(clknet_leaf_0_pclk));
 BUF_X4 clkbuf_leaf_1_pclk (.A(clknet_2_0__leaf_pclk),
    .Z(clknet_leaf_1_pclk));
 BUF_X4 clkbuf_leaf_2_pclk (.A(clknet_2_0__leaf_pclk),
    .Z(clknet_leaf_2_pclk));
 BUF_X4 clkbuf_leaf_3_pclk (.A(clknet_2_1__leaf_pclk),
    .Z(clknet_leaf_3_pclk));
 BUF_X4 clkbuf_leaf_4_pclk (.A(clknet_2_1__leaf_pclk),
    .Z(clknet_leaf_4_pclk));
 BUF_X4 clkbuf_leaf_5_pclk (.A(clknet_2_1__leaf_pclk),
    .Z(clknet_leaf_5_pclk));
 BUF_X4 clkbuf_leaf_6_pclk (.A(clknet_2_1__leaf_pclk),
    .Z(clknet_leaf_6_pclk));
 BUF_X4 clkbuf_leaf_7_pclk (.A(clknet_2_1__leaf_pclk),
    .Z(clknet_leaf_7_pclk));
 BUF_X4 clkbuf_leaf_8_pclk (.A(clknet_2_1__leaf_pclk),
    .Z(clknet_leaf_8_pclk));
 BUF_X4 clkbuf_leaf_9_pclk (.A(clknet_2_1__leaf_pclk),
    .Z(clknet_leaf_9_pclk));
 BUF_X4 clkbuf_leaf_10_pclk (.A(clknet_2_1__leaf_pclk),
    .Z(clknet_leaf_10_pclk));
 BUF_X4 clkbuf_leaf_11_pclk (.A(clknet_2_1__leaf_pclk),
    .Z(clknet_leaf_11_pclk));
 BUF_X4 clkbuf_leaf_12_pclk (.A(clknet_2_3__leaf_pclk),
    .Z(clknet_leaf_12_pclk));
 BUF_X4 clkbuf_leaf_13_pclk (.A(clknet_2_3__leaf_pclk),
    .Z(clknet_leaf_13_pclk));
 BUF_X4 clkbuf_leaf_14_pclk (.A(clknet_2_3__leaf_pclk),
    .Z(clknet_leaf_14_pclk));
 BUF_X4 clkbuf_leaf_15_pclk (.A(clknet_2_3__leaf_pclk),
    .Z(clknet_leaf_15_pclk));
 BUF_X4 clkbuf_leaf_16_pclk (.A(clknet_2_3__leaf_pclk),
    .Z(clknet_leaf_16_pclk));
 BUF_X4 clkbuf_leaf_17_pclk (.A(clknet_2_3__leaf_pclk),
    .Z(clknet_leaf_17_pclk));
 BUF_X4 clkbuf_leaf_18_pclk (.A(clknet_2_3__leaf_pclk),
    .Z(clknet_leaf_18_pclk));
 BUF_X4 clkbuf_leaf_19_pclk (.A(clknet_2_3__leaf_pclk),
    .Z(clknet_leaf_19_pclk));
 BUF_X4 clkbuf_leaf_20_pclk (.A(clknet_2_3__leaf_pclk),
    .Z(clknet_leaf_20_pclk));
 BUF_X4 clkbuf_leaf_21_pclk (.A(clknet_2_2__leaf_pclk),
    .Z(clknet_leaf_21_pclk));
 BUF_X4 clkbuf_leaf_22_pclk (.A(clknet_2_2__leaf_pclk),
    .Z(clknet_leaf_22_pclk));
 BUF_X4 clkbuf_leaf_23_pclk (.A(clknet_2_2__leaf_pclk),
    .Z(clknet_leaf_23_pclk));
 BUF_X4 clkbuf_leaf_24_pclk (.A(clknet_2_2__leaf_pclk),
    .Z(clknet_leaf_24_pclk));
 BUF_X4 clkbuf_leaf_25_pclk (.A(clknet_2_2__leaf_pclk),
    .Z(clknet_leaf_25_pclk));
 BUF_X4 clkbuf_leaf_26_pclk (.A(clknet_2_2__leaf_pclk),
    .Z(clknet_leaf_26_pclk));
 BUF_X4 clkbuf_leaf_27_pclk (.A(clknet_2_2__leaf_pclk),
    .Z(clknet_leaf_27_pclk));
 BUF_X4 clkbuf_leaf_28_pclk (.A(clknet_2_2__leaf_pclk),
    .Z(clknet_leaf_28_pclk));
 BUF_X4 clkbuf_leaf_29_pclk (.A(clknet_2_2__leaf_pclk),
    .Z(clknet_leaf_29_pclk));
 BUF_X4 clkbuf_leaf_30_pclk (.A(clknet_2_0__leaf_pclk),
    .Z(clknet_leaf_30_pclk));
 BUF_X4 clkbuf_leaf_31_pclk (.A(clknet_2_0__leaf_pclk),
    .Z(clknet_leaf_31_pclk));
 BUF_X4 clkbuf_leaf_32_pclk (.A(clknet_2_0__leaf_pclk),
    .Z(clknet_leaf_32_pclk));
 BUF_X4 clkbuf_leaf_33_pclk (.A(clknet_2_0__leaf_pclk),
    .Z(clknet_leaf_33_pclk));
 BUF_X4 clkbuf_leaf_34_pclk (.A(clknet_2_0__leaf_pclk),
    .Z(clknet_leaf_34_pclk));
 BUF_X4 clkbuf_leaf_35_pclk (.A(clknet_2_0__leaf_pclk),
    .Z(clknet_leaf_35_pclk));
 BUF_X4 clkbuf_0_pclk (.A(pclk),
    .Z(clknet_0_pclk));
 BUF_X4 clkbuf_2_0__f_pclk (.A(clknet_0_pclk),
    .Z(clknet_2_0__leaf_pclk));
 BUF_X4 clkbuf_2_1__f_pclk (.A(clknet_0_pclk),
    .Z(clknet_2_1__leaf_pclk));
 BUF_X4 clkbuf_2_2__f_pclk (.A(clknet_0_pclk),
    .Z(clknet_2_2__leaf_pclk));
 BUF_X4 clkbuf_2_3__f_pclk (.A(clknet_0_pclk),
    .Z(clknet_2_3__leaf_pclk));
 INV_X1 clkload0 (.A(clknet_leaf_0_pclk));
 INV_X1 clkload1 (.A(clknet_leaf_2_pclk));
 INV_X1 clkload2 (.A(clknet_leaf_30_pclk));
 INV_X1 clkload3 (.A(clknet_leaf_31_pclk));
 INV_X1 clkload4 (.A(clknet_leaf_32_pclk));
 INV_X1 clkload5 (.A(clknet_leaf_33_pclk));
 INV_X1 clkload6 (.A(clknet_leaf_34_pclk));
 INV_X16 clkload7 (.A(clknet_leaf_35_pclk));
 INV_X1 clkload8 (.A(clknet_leaf_3_pclk));
 INV_X1 clkload9 (.A(clknet_leaf_4_pclk));
 INV_X1 clkload10 (.A(clknet_leaf_6_pclk));
 INV_X1 clkload11 (.A(clknet_leaf_7_pclk));
 INV_X1 clkload12 (.A(clknet_leaf_8_pclk));
 INV_X1 clkload13 (.A(clknet_leaf_9_pclk));
 INV_X1 clkload14 (.A(clknet_leaf_10_pclk));
 INV_X1 clkload15 (.A(clknet_leaf_11_pclk));
 INV_X1 clkload16 (.A(clknet_leaf_21_pclk));
 INV_X1 clkload17 (.A(clknet_leaf_22_pclk));
 INV_X1 clkload18 (.A(clknet_leaf_23_pclk));
 INV_X1 clkload19 (.A(clknet_leaf_24_pclk));
 INV_X1 clkload20 (.A(clknet_leaf_26_pclk));
 INV_X1 clkload21 (.A(clknet_leaf_27_pclk));
 INV_X1 clkload22 (.A(clknet_leaf_28_pclk));
 INV_X1 clkload23 (.A(clknet_leaf_29_pclk));
 INV_X1 clkload24 (.A(clknet_leaf_12_pclk));
 INV_X1 clkload25 (.A(clknet_leaf_13_pclk));
 INV_X1 clkload26 (.A(clknet_leaf_14_pclk));
 INV_X1 clkload27 (.A(clknet_leaf_15_pclk));
 INV_X1 clkload28 (.A(clknet_leaf_16_pclk));
 INV_X1 clkload29 (.A(clknet_leaf_17_pclk));
 INV_X1 clkload30 (.A(clknet_leaf_19_pclk));
 INV_X1 clkload31 (.A(clknet_leaf_20_pclk));
 BUF_X1 hold71 (.A(_0000_),
    .Z(net71));
 assign temp[0] = prdata[0];
 assign temp[10] = prdata[10];
 assign temp[11] = prdata[11];
 assign temp[12] = prdata[12];
 assign temp[13] = prdata[13];
 assign temp[14] = prdata[14];
 assign temp[15] = prdata[15];
 assign temp[16] = prdata[16];
 assign temp[17] = prdata[17];
 assign temp[18] = prdata[18];
 assign temp[19] = prdata[19];
 assign temp[1] = prdata[1];
 assign temp[20] = prdata[20];
 assign temp[21] = prdata[21];
 assign temp[22] = prdata[22];
 assign temp[23] = prdata[23];
 assign temp[24] = prdata[24];
 assign temp[25] = prdata[25];
 assign temp[26] = prdata[26];
 assign temp[27] = prdata[27];
 assign temp[28] = prdata[28];
 assign temp[29] = prdata[29];
 assign temp[2] = prdata[2];
 assign temp[30] = prdata[30];
 assign temp[31] = prdata[31];
 assign temp[3] = prdata[3];
 assign temp[4] = prdata[4];
 assign temp[5] = prdata[5];
 assign temp[6] = prdata[6];
 assign temp[7] = prdata[7];
 assign temp[8] = prdata[8];
 assign temp[9] = prdata[9];
endmodule
