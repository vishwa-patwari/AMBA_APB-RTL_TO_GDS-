module apb_memory_tb;
  reg pclk;
  reg prst_n;
  reg pselx;
  reg penable;
  reg pwrite;
  reg [31:0] pwdata;
  reg [31:0] paddr;

  wire pready;
  wire pslverr;
  wire [31:0] prdata;
  wire [31:0] temp;

  // Store last written addr for readback
  reg [31:0] last_addr;

  // DUT Instance
  apb_slave_memory dut (
    .pclk(pclk), .prst_n(prst_n), .paddr(paddr),
    .pselx(pselx), .penable(penable), .pwrite(pwrite),
    .pwdata(pwdata), .pready(pready), .pslverr(pslverr),
    .prdata(prdata), .temp(temp)
  );

  ////// Clock generation ////// 
  initial pclk = 1;
  always #10 pclk = ~pclk;

  ////// Reset and initialization ///////
  task reset_and_initialization;
    begin
      #5 prst_n = 0;
      @(posedge pclk);
      prst_n = 1;
      pselx  = 0;
      penable = 0;
      pwrite = 0;
      pwdata = 0;
      paddr  = 0;
    end
  endtask

  ////// Write transfer ////// 
  task write_transfer;
    begin
      pselx  = 1;
      pwrite = 1;
      pwdata = $random;       // random data
     paddr  = $urandom_range(0, 31);  // valid range 0–31
      last_addr = paddr;      // save addr for readback

      @(posedge pclk);
      penable = 1;

      wait (pready == 1);

      @(posedge pclk);
      penable = 0;

      $strobe("Writing data into memory: data = %0h, address = %0d", pwdata, paddr);
    end
  endtask

  ////// Read transfer ////// 
  task read_transfer;
    begin
      pselx  = 1;
      pwrite = 0;
      paddr  = last_addr;   // read from same addr as last write

      @(posedge pclk);
      penable = 1;

      wait (pready == 1);

      @(posedge pclk);
      pselx  = 0;
      pwrite = 0;
      penable = 0;

      $strobe("Reading data from memory: data = %0h, address = %0d", prdata, paddr);
    end
  endtask

  ////// Read-Write transaction ////// 
  task read_write_transfer;
    begin
      repeat (5) begin      // try 5 random transactions
        write_transfer;
        read_transfer;
      end
    end
  endtask

  //// Initial simulation //// 
  initial begin
    reset_and_initialization;
    read_write_transfer;
    #100 $finish;
  end

  initial begin
    $dumpfile("dump.vcd");
    $dumpvars(0, apb_memory_tb);
  end
endmodule
